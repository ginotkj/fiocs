Analisis Inyeccion VA=3v Afalla=5mA

**** 04/11/10 20:49:07 ******* PSpice 16.0.0 (July 2006) ****** ID# 0 ********

 ** Profile: "PRUEBA-transient"  [ D:\Documents\TESIS\fiocs\Design\I-FLASH-01\OrCAD\I-FLASH-6BITS\i-flash-6bits-pspicefiles\prueba\tr


 ****     CIRCUIT DESCRIPTION


******************************************************************************




** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB D:\Documents\TESIS\fiocs\Design\I-FLASH-01\OrCAD\I-FLASH-6BITS\i-flash-6bits-PSpiceFiles\i-flash-6bits.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.0\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 15n 0 1p 
.OPTIONS NODE
.OPTIONS ITL1= 300
.OPTIONS ITL2= 100
.PROBE
*.INC "..\PRUEBA.net" 



**** INCLUDING PRUEBA.net ****
* source I-FLASH-6BITS
R_R6         LSB N116990  100k  
R_R7         N-MSB N116990  100k  
V_Clock         N116976 0  
+PULSE 0 3 .4u 0.05u 0.05u .4u 1u
R_R8         N-5SB N116990  100k  
M_CONV_FLASH_C38_M4         CONV_FLASH_C38_ND+ CONV_FLASH_C38_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C38_M5         CONV_FLASH_C38_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C38_M6         Q38 CONV_FLASH_C38_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C38_M7         Q38 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C38_M1         CONV_FLASH_C38_ND- N117007 CONV_FLASH_C38_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C38_M2         CONV_FLASH_C38_ND+ CONV_N117508
+  CONV_FLASH_C38_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C38_M3         CONV_FLASH_C38_ND- CONV_FLASH_C38_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C5_M4         CONV_FLASH_C5_ND+ CONV_FLASH_C5_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C5_M5         CONV_FLASH_C5_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C5_M6         Q5 CONV_FLASH_C5_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C5_M7         Q5 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C5_M1         CONV_FLASH_C5_ND- N117007 CONV_FLASH_C5_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C5_M2         CONV_FLASH_C5_ND+ CONV_N117574 CONV_FLASH_C5_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C5_M3         CONV_FLASH_C5_ND- CONV_FLASH_C5_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C25_M4         CONV_FLASH_C25_ND+ CONV_FLASH_C25_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C25_M5         CONV_FLASH_C25_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C25_M6         Q25 CONV_FLASH_C25_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C25_M7         Q25 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C25_M1         CONV_FLASH_C25_ND- N117007 CONV_FLASH_C25_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C25_M2         CONV_FLASH_C25_ND+ CONV_N117534
+  CONV_FLASH_C25_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C25_M3         CONV_FLASH_C25_ND- CONV_FLASH_C25_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C31_M4         CONV_FLASH_C31_ND+ CONV_FLASH_C31_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C31_M5         CONV_FLASH_C31_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C31_M6         Q31 CONV_FLASH_C31_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C31_M7         Q31 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C31_M1         CONV_FLASH_C31_ND- N117007 CONV_FLASH_C31_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C31_M2         CONV_FLASH_C31_ND+ CONV_N117522
+  CONV_FLASH_C31_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C31_M3         CONV_FLASH_C31_ND- CONV_FLASH_C31_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C8_M4         CONV_FLASH_C8_ND+ CONV_FLASH_C8_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C8_M5         CONV_FLASH_C8_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C8_M6         Q8 CONV_FLASH_C8_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C8_M7         Q8 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C8_M1         CONV_FLASH_C8_ND- N117007 CONV_FLASH_C8_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C8_M2         CONV_FLASH_C8_ND+ CONV_N117576 CONV_FLASH_C8_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C8_M3         CONV_FLASH_C8_ND- CONV_FLASH_C8_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C19_M4         CONV_FLASH_C19_ND+ CONV_FLASH_C19_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C19_M5         CONV_FLASH_C19_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C19_M6         Q19 CONV_FLASH_C19_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C19_M7         Q19 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C19_M1         CONV_FLASH_C19_ND- N117007 CONV_FLASH_C19_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C19_M2         CONV_FLASH_C19_ND+ CONV_N117546
+  CONV_FLASH_C19_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C19_M3         CONV_FLASH_C19_ND- CONV_FLASH_C19_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C2_M4         CONV_FLASH_C2_ND+ CONV_FLASH_C2_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C2_M5         CONV_FLASH_C2_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C2_M6         Q2 CONV_FLASH_C2_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C2_M7         Q2 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C2_M1         CONV_FLASH_C2_ND- N117007 CONV_FLASH_C2_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C2_M2         CONV_FLASH_C2_ND+ CONV_N117564 CONV_FLASH_C2_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C2_M3         CONV_FLASH_C2_ND- CONV_FLASH_C2_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C46_M4         CONV_FLASH_C46_ND+ CONV_FLASH_C46_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C46_M5         CONV_FLASH_C46_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C46_M6         Q46 CONV_FLASH_C46_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C46_M7         Q46 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C46_M1         CONV_FLASH_C46_ND- N117007 CONV_FLASH_C46_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C46_M2         CONV_FLASH_C46_ND+ CONV_N117494
+  CONV_FLASH_C46_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C46_M3         CONV_FLASH_C46_ND- CONV_FLASH_C46_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C47_M4         CONV_FLASH_C47_ND+ CONV_FLASH_C47_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C47_M5         CONV_FLASH_C47_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C47_M6         Q47 CONV_FLASH_C47_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C47_M7         Q47 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C47_M1         CONV_FLASH_C47_ND- N117007 CONV_FLASH_C47_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C47_M2         CONV_FLASH_C47_ND+ CONV_N117496
+  CONV_FLASH_C47_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C47_M3         CONV_FLASH_C47_ND- CONV_FLASH_C47_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C60_M4         CONV_FLASH_C60_ND+ CONV_FLASH_C60_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C60_M5         CONV_FLASH_C60_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C60_M6         Q60 CONV_FLASH_C60_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C60_M7         Q60 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C60_M1         CONV_FLASH_C60_ND- N117007 CONV_FLASH_C60_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C60_M2         CONV_FLASH_C60_ND+ CONV_N119887
+  CONV_FLASH_C60_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C60_M3         CONV_FLASH_C60_ND- CONV_FLASH_C60_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C45_M4         CONV_FLASH_C45_ND+ CONV_FLASH_C45_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C45_M5         CONV_FLASH_C45_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C45_M6         Q45 CONV_FLASH_C45_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C45_M7         Q45 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C45_M1         CONV_FLASH_C45_ND- N117007 CONV_FLASH_C45_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C45_M2         CONV_FLASH_C45_ND+ CONV_N117492
+  CONV_FLASH_C45_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C45_M3         CONV_FLASH_C45_ND- CONV_FLASH_C45_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C54_M4         CONV_FLASH_C54_ND+ CONV_FLASH_C54_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C54_M5         CONV_FLASH_C54_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C54_M6         Q54 CONV_FLASH_C54_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C54_M7         Q54 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C54_M1         CONV_FLASH_C54_ND- N117007 CONV_FLASH_C54_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C54_M2         CONV_FLASH_C54_ND+ CONV_N119899
+  CONV_FLASH_C54_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C54_M3         CONV_FLASH_C54_ND- CONV_FLASH_C54_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C34_M4         CONV_FLASH_C34_ND+ CONV_FLASH_C34_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C34_M5         CONV_FLASH_C34_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C34_M6         Q34 CONV_FLASH_C34_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C34_M7         Q34 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C34_M1         CONV_FLASH_C34_ND- N117007 CONV_FLASH_C34_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C34_M2         CONV_FLASH_C34_ND+ CONV_N117516
+  CONV_FLASH_C34_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C34_M3         CONV_FLASH_C34_ND- CONV_FLASH_C34_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C26_M4         CONV_FLASH_C26_ND+ CONV_FLASH_C26_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C26_M5         CONV_FLASH_C26_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C26_M6         Q26 CONV_FLASH_C26_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C26_M7         Q26 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C26_M1         CONV_FLASH_C26_ND- N117007 CONV_FLASH_C26_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C26_M2         CONV_FLASH_C26_ND+ CONV_N117536
+  CONV_FLASH_C26_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C26_M3         CONV_FLASH_C26_ND- CONV_FLASH_C26_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C48_M4         CONV_FLASH_C48_ND+ CONV_FLASH_C48_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C48_M5         CONV_FLASH_C48_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C48_M6         Q48 CONV_FLASH_C48_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C48_M7         Q48 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C48_M1         CONV_FLASH_C48_ND- N117007 CONV_FLASH_C48_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C48_M2         CONV_FLASH_C48_ND+ CONV_N117498
+  CONV_FLASH_C48_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C48_M3         CONV_FLASH_C48_ND- CONV_FLASH_C48_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C44_M4         CONV_FLASH_C44_ND+ CONV_FLASH_C44_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C44_M5         CONV_FLASH_C44_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C44_M6         Q44 CONV_FLASH_C44_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C44_M7         Q44 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C44_M1         CONV_FLASH_C44_ND- N117007 CONV_FLASH_C44_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C44_M2         CONV_FLASH_C44_ND+ CONV_N117490
+  CONV_FLASH_C44_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C44_M3         CONV_FLASH_C44_ND- CONV_FLASH_C44_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C7_M4         CONV_FLASH_C7_ND+ CONV_FLASH_C7_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C7_M5         CONV_FLASH_C7_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C7_M6         Q7 CONV_FLASH_C7_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C7_M7         Q7 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C7_M1         CONV_FLASH_C7_ND- N117007 CONV_FLASH_C7_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C7_M2         CONV_FLASH_C7_ND+ CONV_N117570 CONV_FLASH_C7_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C7_M3         CONV_FLASH_C7_ND- CONV_FLASH_C7_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C18_M4         CONV_FLASH_C18_ND+ CONV_FLASH_C18_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C18_M5         CONV_FLASH_C18_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C18_M6         Q18 CONV_FLASH_C18_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C18_M7         Q18 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C18_M1         CONV_FLASH_C18_ND- N117007 CONV_FLASH_C18_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C18_M2         CONV_FLASH_C18_ND+ CONV_N117548
+  CONV_FLASH_C18_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C18_M3         CONV_FLASH_C18_ND- CONV_FLASH_C18_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_FFD6_NAND6_M5         CONV_FLASH_FFD6_N62152 CONV_FLASH_FFD6_Y
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND6_M6         CONV_FLASH_FFD6_N62152 CONV_FLASH_FFD6_Y
+  CONV_FLASH_FFD6_NAND6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND6_M2         CONV_FLASH_FFD6_NAND6_ND2 CONV_FLASH_D-MSB 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND6_M4         CONV_FLASH_FFD6_N62152 CONV_FLASH_D-MSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND1_M2         CONV_FLASH_FFD6_NAND1_ND2 N116976
+  CONV_FLASH_FFD6_NAND1_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND1_M3         CONV_FLASH_FFD6_Y CONV_FLASH_FFD6_X N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND1_M6         CONV_FLASH_FFD6_NAND1_ND3
+  CONV_FLASH_FFD6_N62152 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND1_M4         CONV_FLASH_FFD6_Y N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND1_M1         CONV_FLASH_FFD6_Y CONV_FLASH_FFD6_X
+  CONV_FLASH_FFD6_NAND1_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND1_M5         CONV_FLASH_FFD6_Y CONV_FLASH_FFD6_N62152
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND2_M5         CONV_FLASH_FFD6_N62128
+  CONV_FLASH_FFD6_N62152 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND2_M6         CONV_FLASH_FFD6_N62128
+  CONV_FLASH_FFD6_N62152 CONV_FLASH_FFD6_NAND2_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND2_M2         CONV_FLASH_FFD6_NAND2_ND2 CONV_FLASH_FFD6_X
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND2_M4         CONV_FLASH_FFD6_N62128 CONV_FLASH_FFD6_X
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND3_M5         CONV_FLASH_FFD6_X CONV_FLASH_FFD6_N62128
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND3_M6         CONV_FLASH_FFD6_X CONV_FLASH_FFD6_N62128
+  CONV_FLASH_FFD6_NAND3_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND3_M2         CONV_FLASH_FFD6_NAND3_ND2 N116976 0 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND3_M4         CONV_FLASH_FFD6_X N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND4_M5         MSB CONV_FLASH_FFD6_X N116990 N116990 CMOSP 
+  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND4_M6         MSB CONV_FLASH_FFD6_X
+  CONV_FLASH_FFD6_NAND4_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND4_M2         CONV_FLASH_FFD6_NAND4_ND2 N-MSB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND4_M4         MSB N-MSB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND5_M5         N-MSB MSB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD6_NAND5_M6         N-MSB MSB CONV_FLASH_FFD6_NAND5_ND2 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND5_M2         CONV_FLASH_FFD6_NAND5_ND2 CONV_FLASH_FFD6_Y
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD6_NAND5_M4         N-MSB CONV_FLASH_FFD6_Y N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_C4_M4         CONV_FLASH_C4_ND+ CONV_FLASH_C4_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C4_M5         CONV_FLASH_C4_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C4_M6         Q4 CONV_FLASH_C4_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C4_M7         Q4 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C4_M1         CONV_FLASH_C4_ND- N117007 CONV_FLASH_C4_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C4_M2         CONV_FLASH_C4_ND+ CONV_N117566 CONV_FLASH_C4_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C4_M3         CONV_FLASH_C4_ND- CONV_FLASH_C4_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C49_M4         CONV_FLASH_C49_ND+ CONV_FLASH_C49_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C49_M5         CONV_FLASH_C49_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C49_M6         Q49 CONV_FLASH_C49_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C49_M7         Q49 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C49_M1         CONV_FLASH_C49_ND- N117007 CONV_FLASH_C49_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C49_M2         CONV_FLASH_C49_ND+ CONV_N117500
+  CONV_FLASH_C49_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C49_M3         CONV_FLASH_C49_ND- CONV_FLASH_C49_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C43_M4         CONV_FLASH_C43_ND+ CONV_FLASH_C43_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C43_M5         CONV_FLASH_C43_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C43_M6         Q43 CONV_FLASH_C43_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C43_M7         Q43 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C43_M1         CONV_FLASH_C43_ND- N117007 CONV_FLASH_C43_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C43_M2         CONV_FLASH_C43_ND+ CONV_N117488
+  CONV_FLASH_C43_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C43_M3         CONV_FLASH_C43_ND- CONV_FLASH_C43_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C37_M4         CONV_FLASH_C37_ND+ CONV_FLASH_C37_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C37_M5         CONV_FLASH_C37_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C37_M6         Q37 CONV_FLASH_C37_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C37_M7         Q37 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C37_M1         CONV_FLASH_C37_ND- N117007 CONV_FLASH_C37_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C37_M2         CONV_FLASH_C37_ND+ CONV_N117510
+  CONV_FLASH_C37_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C37_M3         CONV_FLASH_C37_ND- CONV_FLASH_C37_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C27_M4         CONV_FLASH_C27_ND+ CONV_FLASH_C27_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C27_M5         CONV_FLASH_C27_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C27_M6         Q27 CONV_FLASH_C27_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C27_M7         Q27 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C27_M1         CONV_FLASH_C27_ND- N117007 CONV_FLASH_C27_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C27_M2         CONV_FLASH_C27_ND+ CONV_N117538
+  CONV_FLASH_C27_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C27_M3         CONV_FLASH_C27_ND- CONV_FLASH_C27_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_FFD3_NAND6_M5         CONV_FLASH_FFD3_N62152 CONV_FLASH_FFD3_Y
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND6_M6         CONV_FLASH_FFD3_N62152 CONV_FLASH_FFD3_Y
+  CONV_FLASH_FFD3_NAND6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND6_M2         CONV_FLASH_FFD3_NAND6_ND2 CONV_FLASH_D-3SB 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND6_M4         CONV_FLASH_FFD3_N62152 CONV_FLASH_D-3SB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND1_M2         CONV_FLASH_FFD3_NAND1_ND2 N116976
+  CONV_FLASH_FFD3_NAND1_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND1_M3         CONV_FLASH_FFD3_Y CONV_FLASH_FFD3_X N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND1_M6         CONV_FLASH_FFD3_NAND1_ND3
+  CONV_FLASH_FFD3_N62152 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND1_M4         CONV_FLASH_FFD3_Y N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND1_M1         CONV_FLASH_FFD3_Y CONV_FLASH_FFD3_X
+  CONV_FLASH_FFD3_NAND1_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND1_M5         CONV_FLASH_FFD3_Y CONV_FLASH_FFD3_N62152
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND2_M5         CONV_FLASH_FFD3_N62128
+  CONV_FLASH_FFD3_N62152 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND2_M6         CONV_FLASH_FFD3_N62128
+  CONV_FLASH_FFD3_N62152 CONV_FLASH_FFD3_NAND2_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND2_M2         CONV_FLASH_FFD3_NAND2_ND2 CONV_FLASH_FFD3_X
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND2_M4         CONV_FLASH_FFD3_N62128 CONV_FLASH_FFD3_X
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND3_M5         CONV_FLASH_FFD3_X CONV_FLASH_FFD3_N62128
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND3_M6         CONV_FLASH_FFD3_X CONV_FLASH_FFD3_N62128
+  CONV_FLASH_FFD3_NAND3_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND3_M2         CONV_FLASH_FFD3_NAND3_ND2 N116976 0 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND3_M4         CONV_FLASH_FFD3_X N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND4_M5         3SB CONV_FLASH_FFD3_X N116990 N116990 CMOSP 
+  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND4_M6         3SB CONV_FLASH_FFD3_X
+  CONV_FLASH_FFD3_NAND4_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND4_M2         CONV_FLASH_FFD3_NAND4_ND2 N-3SB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND4_M4         3SB N-3SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND5_M5         N-3SB 3SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD3_NAND5_M6         N-3SB 3SB CONV_FLASH_FFD3_NAND5_ND2 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND5_M2         CONV_FLASH_FFD3_NAND5_ND2 CONV_FLASH_FFD3_Y
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD3_NAND5_M4         N-3SB CONV_FLASH_FFD3_Y N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_C32_M4         CONV_FLASH_C32_ND+ CONV_FLASH_C32_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C32_M5         CONV_FLASH_C32_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C32_M6         CONV_FLASH_D-MSB CONV_FLASH_C32_ND+ N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C32_M7         CONV_FLASH_D-MSB N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C32_M1         CONV_FLASH_C32_ND- N117007 CONV_FLASH_C32_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C32_M2         CONV_FLASH_C32_ND+ CONV_N117520
+  CONV_FLASH_C32_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C32_M3         CONV_FLASH_C32_ND- CONV_FLASH_C32_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C58_M4         CONV_FLASH_C58_ND+ CONV_FLASH_C58_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C58_M5         CONV_FLASH_C58_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C58_M6         Q58 CONV_FLASH_C58_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C58_M7         Q58 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C58_M1         CONV_FLASH_C58_ND- N117007 CONV_FLASH_C58_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C58_M2         CONV_FLASH_C58_ND+ CONV_N119891
+  CONV_FLASH_C58_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C58_M3         CONV_FLASH_C58_ND- CONV_FLASH_C58_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C17_M4         CONV_FLASH_C17_ND+ CONV_FLASH_C17_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C17_M5         CONV_FLASH_C17_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C17_M6         Q17 CONV_FLASH_C17_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C17_M7         Q17 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C17_M1         CONV_FLASH_C17_ND- N117007 CONV_FLASH_C17_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C17_M2         CONV_FLASH_C17_ND+ CONV_N117550
+  CONV_FLASH_C17_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C17_M3         CONV_FLASH_C17_ND- CONV_FLASH_C17_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C42_M4         CONV_FLASH_C42_ND+ CONV_FLASH_C42_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C42_M5         CONV_FLASH_C42_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C42_M6         Q42 CONV_FLASH_C42_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C42_M7         Q42 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C42_M1         CONV_FLASH_C42_ND- N117007 CONV_FLASH_C42_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C42_M2         CONV_FLASH_C42_ND+ CONV_N117486
+  CONV_FLASH_C42_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C42_M3         CONV_FLASH_C42_ND- CONV_FLASH_C42_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C50_M4         CONV_FLASH_C50_ND+ CONV_FLASH_C50_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C50_M5         CONV_FLASH_C50_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C50_M6         Q50 CONV_FLASH_C50_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C50_M7         Q50 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C50_M1         CONV_FLASH_C50_ND- N117007 CONV_FLASH_C50_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C50_M2         CONV_FLASH_C50_ND+ CONV_N119903
+  CONV_FLASH_C50_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C50_M3         CONV_FLASH_C50_ND- CONV_FLASH_C50_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C55_M4         CONV_FLASH_C55_ND+ CONV_FLASH_C55_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C55_M5         CONV_FLASH_C55_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C55_M6         Q55 CONV_FLASH_C55_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C55_M7         Q55 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C55_M1         CONV_FLASH_C55_ND- N117007 CONV_FLASH_C55_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C55_M2         CONV_FLASH_C55_ND+ CONV_N119897
+  CONV_FLASH_C55_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C55_M3         CONV_FLASH_C55_ND- CONV_FLASH_C55_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C3_M4         CONV_FLASH_C3_ND+ CONV_FLASH_C3_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C3_M5         CONV_FLASH_C3_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C3_M6         Q3 CONV_FLASH_C3_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C3_M7         Q3 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C3_M1         CONV_FLASH_C3_ND- N117007 CONV_FLASH_C3_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C3_M2         CONV_FLASH_C3_ND+ CONV_N117568 CONV_FLASH_C3_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C3_M3         CONV_FLASH_C3_ND- CONV_FLASH_C3_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C28_M4         CONV_FLASH_C28_ND+ CONV_FLASH_C28_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C28_M5         CONV_FLASH_C28_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C28_M6         Q28 CONV_FLASH_C28_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C28_M7         Q28 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C28_M1         CONV_FLASH_C28_ND- N117007 CONV_FLASH_C28_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C28_M2         CONV_FLASH_C28_ND+ CONV_N117540
+  CONV_FLASH_C28_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C28_M3         CONV_FLASH_C28_ND- CONV_FLASH_C28_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C63_M4         CONV_FLASH_C63_ND+ CONV_FLASH_C63_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C63_M5         CONV_FLASH_C63_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C63_M6         Q63 CONV_FLASH_C63_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C63_M7         Q63 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C63_M1         CONV_FLASH_C63_ND- N117007 CONV_FLASH_C63_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C63_M2         CONV_FLASH_C63_ND+ CONV_N119881
+  CONV_FLASH_C63_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C63_M3         CONV_FLASH_C63_ND- CONV_FLASH_C63_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C41_M4         CONV_FLASH_C41_ND+ CONV_FLASH_C41_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C41_M5         CONV_FLASH_C41_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C41_M6         Q41 CONV_FLASH_C41_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C41_M7         Q41 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C41_M1         CONV_FLASH_C41_ND- N117007 CONV_FLASH_C41_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C41_M2         CONV_FLASH_C41_ND+ CONV_N117502
+  CONV_FLASH_C41_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C41_M3         CONV_FLASH_C41_ND- CONV_FLASH_C41_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C33_M4         CONV_FLASH_C33_ND+ CONV_FLASH_C33_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C33_M5         CONV_FLASH_C33_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C33_M6         Q33 CONV_FLASH_C33_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C33_M7         Q33 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C33_M1         CONV_FLASH_C33_ND- N117007 CONV_FLASH_C33_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C33_M2         CONV_FLASH_C33_ND+ CONV_N117518
+  CONV_FLASH_C33_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C33_M3         CONV_FLASH_C33_ND- CONV_FLASH_C33_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C51_M4         CONV_FLASH_C51_ND+ CONV_FLASH_C51_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C51_M5         CONV_FLASH_C51_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C51_M6         Q51 CONV_FLASH_C51_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C51_M7         Q51 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C51_M1         CONV_FLASH_C51_ND- N117007 CONV_FLASH_C51_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C51_M2         CONV_FLASH_C51_ND+ CONV_N119905
+  CONV_FLASH_C51_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C51_M3         CONV_FLASH_C51_ND- CONV_FLASH_C51_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C36_M4         CONV_FLASH_C36_ND+ CONV_FLASH_C36_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C36_M5         CONV_FLASH_C36_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C36_M6         Q36 CONV_FLASH_C36_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C36_M7         Q36 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C36_M1         CONV_FLASH_C36_ND- N117007 CONV_FLASH_C36_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C36_M2         CONV_FLASH_C36_ND+ CONV_N117512
+  CONV_FLASH_C36_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C36_M3         CONV_FLASH_C36_ND- CONV_FLASH_C36_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C61_M4         CONV_FLASH_C61_ND+ CONV_FLASH_C61_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C61_M5         CONV_FLASH_C61_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C61_M6         Q61 CONV_FLASH_C61_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C61_M7         Q61 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C61_M1         CONV_FLASH_C61_ND- N117007 CONV_FLASH_C61_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C61_M2         CONV_FLASH_C61_ND+ CONV_N119885
+  CONV_FLASH_C61_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C61_M3         CONV_FLASH_C61_ND- CONV_FLASH_C61_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_FFD4_NAND6_M5         CONV_FLASH_FFD4_N62152 CONV_FLASH_FFD4_Y
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND6_M6         CONV_FLASH_FFD4_N62152 CONV_FLASH_FFD4_Y
+  CONV_FLASH_FFD4_NAND6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND6_M2         CONV_FLASH_FFD4_NAND6_ND2 CONV_FLASH_D-4SB 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND6_M4         CONV_FLASH_FFD4_N62152 CONV_FLASH_D-4SB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND1_M2         CONV_FLASH_FFD4_NAND1_ND2 N116976
+  CONV_FLASH_FFD4_NAND1_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND1_M3         CONV_FLASH_FFD4_Y CONV_FLASH_FFD4_X N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND1_M6         CONV_FLASH_FFD4_NAND1_ND3
+  CONV_FLASH_FFD4_N62152 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND1_M4         CONV_FLASH_FFD4_Y N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND1_M1         CONV_FLASH_FFD4_Y CONV_FLASH_FFD4_X
+  CONV_FLASH_FFD4_NAND1_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND1_M5         CONV_FLASH_FFD4_Y CONV_FLASH_FFD4_N62152
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND2_M5         CONV_FLASH_FFD4_N62128
+  CONV_FLASH_FFD4_N62152 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND2_M6         CONV_FLASH_FFD4_N62128
+  CONV_FLASH_FFD4_N62152 CONV_FLASH_FFD4_NAND2_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND2_M2         CONV_FLASH_FFD4_NAND2_ND2 CONV_FLASH_FFD4_X
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND2_M4         CONV_FLASH_FFD4_N62128 CONV_FLASH_FFD4_X
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND3_M5         CONV_FLASH_FFD4_X CONV_FLASH_FFD4_N62128
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND3_M6         CONV_FLASH_FFD4_X CONV_FLASH_FFD4_N62128
+  CONV_FLASH_FFD4_NAND3_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND3_M2         CONV_FLASH_FFD4_NAND3_ND2 N116976 0 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND3_M4         CONV_FLASH_FFD4_X N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND4_M5         4SB CONV_FLASH_FFD4_X N116990 N116990 CMOSP 
+  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND4_M6         4SB CONV_FLASH_FFD4_X
+  CONV_FLASH_FFD4_NAND4_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND4_M2         CONV_FLASH_FFD4_NAND4_ND2 N-4SB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND4_M4         4SB N-4SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND5_M5         N-4SB 4SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD4_NAND5_M6         N-4SB 4SB CONV_FLASH_FFD4_NAND5_ND2 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND5_M2         CONV_FLASH_FFD4_NAND5_ND2 CONV_FLASH_FFD4_Y
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD4_NAND5_M4         N-4SB CONV_FLASH_FFD4_Y N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_C29_M4         CONV_FLASH_C29_ND+ CONV_FLASH_C29_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C29_M5         CONV_FLASH_C29_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C29_M6         Q29 CONV_FLASH_C29_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C29_M7         Q29 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C29_M1         CONV_FLASH_C29_ND- N117007 CONV_FLASH_C29_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C29_M2         CONV_FLASH_C29_ND+ CONV_N117542
+  CONV_FLASH_C29_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C29_M3         CONV_FLASH_C29_ND- CONV_FLASH_C29_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C40_M4         CONV_FLASH_C40_ND+ CONV_FLASH_C40_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C40_M5         CONV_FLASH_C40_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C40_M6         Q40 CONV_FLASH_C40_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C40_M7         Q40 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C40_M1         CONV_FLASH_C40_ND- N117007 CONV_FLASH_C40_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C40_M2         CONV_FLASH_C40_ND+ CONV_N117504
+  CONV_FLASH_C40_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C40_M3         CONV_FLASH_C40_ND- CONV_FLASH_C40_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_FFD1_NAND6_M5         CONV_FLASH_FFD1_N62152 CONV_FLASH_FFD1_Y
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND6_M6         CONV_FLASH_FFD1_N62152 CONV_FLASH_FFD1_Y
+  CONV_FLASH_FFD1_NAND6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND6_M2         CONV_FLASH_FFD1_NAND6_ND2 CONV_FLASH_D-LSB 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND6_M4         CONV_FLASH_FFD1_N62152 CONV_FLASH_D-LSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND1_M2         CONV_FLASH_FFD1_NAND1_ND2 N116976
+  CONV_FLASH_FFD1_NAND1_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND1_M3         CONV_FLASH_FFD1_Y CONV_FLASH_FFD1_X N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND1_M6         CONV_FLASH_FFD1_NAND1_ND3
+  CONV_FLASH_FFD1_N62152 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND1_M4         CONV_FLASH_FFD1_Y N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND1_M1         CONV_FLASH_FFD1_Y CONV_FLASH_FFD1_X
+  CONV_FLASH_FFD1_NAND1_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND1_M5         CONV_FLASH_FFD1_Y CONV_FLASH_FFD1_N62152
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND2_M5         CONV_FLASH_FFD1_N62128
+  CONV_FLASH_FFD1_N62152 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND2_M6         CONV_FLASH_FFD1_N62128
+  CONV_FLASH_FFD1_N62152 CONV_FLASH_FFD1_NAND2_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND2_M2         CONV_FLASH_FFD1_NAND2_ND2 CONV_FLASH_FFD1_X
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND2_M4         CONV_FLASH_FFD1_N62128 CONV_FLASH_FFD1_X
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND3_M5         CONV_FLASH_FFD1_X CONV_FLASH_FFD1_N62128
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND3_M6         CONV_FLASH_FFD1_X CONV_FLASH_FFD1_N62128
+  CONV_FLASH_FFD1_NAND3_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND3_M2         CONV_FLASH_FFD1_NAND3_ND2 N116976 0 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND3_M4         CONV_FLASH_FFD1_X N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND4_M5         LSB CONV_FLASH_FFD1_X N116990 N116990 CMOSP 
+  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND4_M6         LSB CONV_FLASH_FFD1_X
+  CONV_FLASH_FFD1_NAND4_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND4_M2         CONV_FLASH_FFD1_NAND4_ND2 N-LSB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND4_M4         LSB N-LSB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND5_M5         N-LSB LSB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD1_NAND5_M6         N-LSB LSB CONV_FLASH_FFD1_NAND5_ND2 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND5_M2         CONV_FLASH_FFD1_NAND5_ND2 CONV_FLASH_FFD1_Y
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD1_NAND5_M4         N-LSB CONV_FLASH_FFD1_Y N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_C56_M4         CONV_FLASH_C56_ND+ CONV_FLASH_C56_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C56_M5         CONV_FLASH_C56_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C56_M6         Q56 CONV_FLASH_C56_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C56_M7         Q56 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C56_M1         CONV_FLASH_C56_ND- N117007 CONV_FLASH_C56_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C56_M2         CONV_FLASH_C56_ND+ CONV_N119895
+  CONV_FLASH_C56_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C56_M3         CONV_FLASH_C56_ND- CONV_FLASH_C56_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C52_M4         CONV_FLASH_C52_ND+ CONV_FLASH_C52_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C52_M5         CONV_FLASH_C52_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C52_M6         Q52 CONV_FLASH_C52_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C52_M7         Q52 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C52_M1         CONV_FLASH_C52_ND- N117007 CONV_FLASH_C52_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C52_M2         CONV_FLASH_C52_ND+ CONV_N119907
+  CONV_FLASH_C52_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C52_M3         CONV_FLASH_C52_ND- CONV_FLASH_C52_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C59_M4         CONV_FLASH_C59_ND+ CONV_FLASH_C59_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C59_M5         CONV_FLASH_C59_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C59_M6         Q59 CONV_FLASH_C59_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C59_M7         Q59 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C59_M1         CONV_FLASH_C59_ND- N117007 CONV_FLASH_C59_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C59_M2         CONV_FLASH_C59_ND+ CONV_N119889
+  CONV_FLASH_C59_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C59_M3         CONV_FLASH_C59_ND- CONV_FLASH_C59_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C13_M4         CONV_FLASH_C13_ND+ CONV_FLASH_C13_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C13_M5         CONV_FLASH_C13_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C13_M6         Q13 CONV_FLASH_C13_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C13_M7         Q13 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C13_M1         CONV_FLASH_C13_ND- N117007 CONV_FLASH_C13_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C13_M2         CONV_FLASH_C13_ND+ CONV_N117558
+  CONV_FLASH_C13_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C13_M3         CONV_FLASH_C13_ND- CONV_FLASH_C13_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C14_M4         CONV_FLASH_C14_ND+ CONV_FLASH_C14_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C14_M5         CONV_FLASH_C14_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C14_M6         Q14 CONV_FLASH_C14_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C14_M7         Q14 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C14_M1         CONV_FLASH_C14_ND- N117007 CONV_FLASH_C14_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C14_M2         CONV_FLASH_C14_ND+ CONV_N117556
+  CONV_FLASH_C14_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C14_M3         CONV_FLASH_C14_ND- CONV_FLASH_C14_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C12_M4         CONV_FLASH_C12_ND+ CONV_FLASH_C12_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C12_M5         CONV_FLASH_C12_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C12_M6         Q12 CONV_FLASH_C12_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C12_M7         Q12 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C12_M1         CONV_FLASH_C12_ND- N117007 CONV_FLASH_C12_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C12_M2         CONV_FLASH_C12_ND+ CONV_N117560
+  CONV_FLASH_C12_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C12_M3         CONV_FLASH_C12_ND- CONV_FLASH_C12_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C30_M4         CONV_FLASH_C30_ND+ CONV_FLASH_C30_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C30_M5         CONV_FLASH_C30_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C30_M6         Q30 CONV_FLASH_C30_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C30_M7         Q30 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C30_M1         CONV_FLASH_C30_ND- N117007 CONV_FLASH_C30_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C30_M2         CONV_FLASH_C30_ND+ CONV_N117544
+  CONV_FLASH_C30_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C30_M3         CONV_FLASH_C30_ND- CONV_FLASH_C30_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C35_M4         CONV_FLASH_C35_ND+ CONV_FLASH_C35_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C35_M5         CONV_FLASH_C35_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C35_M6         Q35 CONV_FLASH_C35_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C35_M7         Q35 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C35_M1         CONV_FLASH_C35_ND- N117007 CONV_FLASH_C35_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C35_M2         CONV_FLASH_C35_ND+ CONV_N117514
+  CONV_FLASH_C35_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C35_M3         CONV_FLASH_C35_ND- CONV_FLASH_C35_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C39_M4         CONV_FLASH_C39_ND+ CONV_FLASH_C39_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C39_M5         CONV_FLASH_C39_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C39_M6         Q39 CONV_FLASH_C39_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C39_M7         Q39 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C39_M1         CONV_FLASH_C39_ND- N117007 CONV_FLASH_C39_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C39_M2         CONV_FLASH_C39_ND+ CONV_N117506
+  CONV_FLASH_C39_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C39_M3         CONV_FLASH_C39_ND- CONV_FLASH_C39_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C15_M4         CONV_FLASH_C15_ND+ CONV_FLASH_C15_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C15_M5         CONV_FLASH_C15_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C15_M6         Q15 CONV_FLASH_C15_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C15_M7         Q15 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C15_M1         CONV_FLASH_C15_ND- N117007 CONV_FLASH_C15_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C15_M2         CONV_FLASH_C15_ND+ CONV_N117554
+  CONV_FLASH_C15_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C15_M3         CONV_FLASH_C15_ND- CONV_FLASH_C15_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C11_M4         CONV_FLASH_C11_ND+ CONV_FLASH_C11_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C11_M5         CONV_FLASH_C11_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C11_M6         Q11 CONV_FLASH_C11_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C11_M7         Q11 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C11_M1         CONV_FLASH_C11_ND- N117007 CONV_FLASH_C11_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C11_M2         CONV_FLASH_C11_ND+ CONV_N117562
+  CONV_FLASH_C11_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C11_M3         CONV_FLASH_C11_ND- CONV_FLASH_C11_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C6_M4         CONV_FLASH_C6_ND+ CONV_FLASH_C6_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C6_M5         CONV_FLASH_C6_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C6_M6         Q6 CONV_FLASH_C6_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C6_M7         Q6 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C6_M1         CONV_FLASH_C6_ND- N117007 CONV_FLASH_C6_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C6_M2         CONV_FLASH_C6_ND+ CONV_N117572 CONV_FLASH_C6_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C6_M3         CONV_FLASH_C6_ND- CONV_FLASH_C6_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C16_M4         CONV_FLASH_C16_ND+ CONV_FLASH_C16_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C16_M5         CONV_FLASH_C16_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C16_M6         Q16 CONV_FLASH_C16_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C16_M7         Q16 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C16_M1         CONV_FLASH_C16_ND- N117007 CONV_FLASH_C16_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C16_M2         CONV_FLASH_C16_ND+ CONV_N117552
+  CONV_FLASH_C16_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C16_M3         CONV_FLASH_C16_ND- CONV_FLASH_C16_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C10_M4         CONV_FLASH_C10_ND+ CONV_FLASH_C10_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C10_M5         CONV_FLASH_C10_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C10_M6         Q10 CONV_FLASH_C10_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C10_M7         Q10 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C10_M1         CONV_FLASH_C10_ND- N117007 CONV_FLASH_C10_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C10_M2         CONV_FLASH_C10_ND+ CONV_N117580
+  CONV_FLASH_C10_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C10_M3         CONV_FLASH_C10_ND- CONV_FLASH_C10_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C53_M4         CONV_FLASH_C53_ND+ CONV_FLASH_C53_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C53_M5         CONV_FLASH_C53_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C53_M6         Q53 CONV_FLASH_C53_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C53_M7         Q53 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C53_M1         CONV_FLASH_C53_ND- N117007 CONV_FLASH_C53_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C53_M2         CONV_FLASH_C53_ND+ CONV_N119901
+  CONV_FLASH_C53_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C53_M3         CONV_FLASH_C53_ND- CONV_FLASH_C53_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_FFD5_NAND6_M5         CONV_FLASH_FFD5_N62152 CONV_FLASH_FFD5_Y
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND6_M6         CONV_FLASH_FFD5_N62152 CONV_FLASH_FFD5_Y
+  CONV_FLASH_FFD5_NAND6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND6_M2         CONV_FLASH_FFD5_NAND6_ND2 CONV_FLASH_D-5SB 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND6_M4         CONV_FLASH_FFD5_N62152 CONV_FLASH_D-5SB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND1_M2         CONV_FLASH_FFD5_NAND1_ND2 N116976
+  CONV_FLASH_FFD5_NAND1_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND1_M3         CONV_FLASH_FFD5_Y CONV_FLASH_FFD5_X N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND1_M6         CONV_FLASH_FFD5_NAND1_ND3
+  CONV_FLASH_FFD5_N62152 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND1_M4         CONV_FLASH_FFD5_Y N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND1_M1         CONV_FLASH_FFD5_Y CONV_FLASH_FFD5_X
+  CONV_FLASH_FFD5_NAND1_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND1_M5         CONV_FLASH_FFD5_Y CONV_FLASH_FFD5_N62152
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND2_M5         CONV_FLASH_FFD5_N62128
+  CONV_FLASH_FFD5_N62152 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND2_M6         CONV_FLASH_FFD5_N62128
+  CONV_FLASH_FFD5_N62152 CONV_FLASH_FFD5_NAND2_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND2_M2         CONV_FLASH_FFD5_NAND2_ND2 CONV_FLASH_FFD5_X
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND2_M4         CONV_FLASH_FFD5_N62128 CONV_FLASH_FFD5_X
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND3_M5         CONV_FLASH_FFD5_X CONV_FLASH_FFD5_N62128
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND3_M6         CONV_FLASH_FFD5_X CONV_FLASH_FFD5_N62128
+  CONV_FLASH_FFD5_NAND3_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND3_M2         CONV_FLASH_FFD5_NAND3_ND2 N116976 0 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND3_M4         CONV_FLASH_FFD5_X N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND4_M5         5SB CONV_FLASH_FFD5_X N116990 N116990 CMOSP 
+  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND4_M6         5SB CONV_FLASH_FFD5_X
+  CONV_FLASH_FFD5_NAND4_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND4_M2         CONV_FLASH_FFD5_NAND4_ND2 N-5SB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND4_M4         5SB N-5SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND5_M5         N-5SB 5SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD5_NAND5_M6         N-5SB 5SB CONV_FLASH_FFD5_NAND5_ND2 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND5_M2         CONV_FLASH_FFD5_NAND5_ND2 CONV_FLASH_FFD5_Y
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD5_NAND5_M4         N-5SB CONV_FLASH_FFD5_Y N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_C22_M4         CONV_FLASH_C22_ND+ CONV_FLASH_C22_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C22_M5         CONV_FLASH_C22_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C22_M6         Q22 CONV_FLASH_C22_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C22_M7         Q22 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C22_M1         CONV_FLASH_C22_ND- N117007 CONV_FLASH_C22_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C22_M2         CONV_FLASH_C22_ND+ CONV_N117528
+  CONV_FLASH_C22_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C22_M3         CONV_FLASH_C22_ND- CONV_FLASH_C22_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C23_M4         CONV_FLASH_C23_ND+ CONV_FLASH_C23_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C23_M5         CONV_FLASH_C23_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C23_M6         Q23 CONV_FLASH_C23_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C23_M7         Q23 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C23_M1         CONV_FLASH_C23_ND- N117007 CONV_FLASH_C23_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C23_M2         CONV_FLASH_C23_ND+ CONV_N117530
+  CONV_FLASH_C23_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C23_M3         CONV_FLASH_C23_ND- CONV_FLASH_C23_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C21_M4         CONV_FLASH_C21_ND+ CONV_FLASH_C21_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C21_M5         CONV_FLASH_C21_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C21_M6         Q21 CONV_FLASH_C21_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C21_M7         Q21 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C21_M1         CONV_FLASH_C21_ND- N117007 CONV_FLASH_C21_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C21_M2         CONV_FLASH_C21_ND+ CONV_N117526
+  CONV_FLASH_C21_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C21_M3         CONV_FLASH_C21_ND- CONV_FLASH_C21_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C1_M4         CONV_FLASH_C1_ND+ CONV_FLASH_C1_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C1_M5         CONV_FLASH_C1_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C1_M6         Q1 CONV_FLASH_C1_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C1_M7         Q1 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C1_M1         CONV_FLASH_C1_ND- N117007 CONV_FLASH_C1_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C1_M2         CONV_FLASH_C1_ND+ CONV_N117582 CONV_FLASH_C1_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C1_M3         CONV_FLASH_C1_ND- CONV_FLASH_C1_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C9_M4         CONV_FLASH_C9_ND+ CONV_FLASH_C9_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C9_M5         CONV_FLASH_C9_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C9_M6         Q9 CONV_FLASH_C9_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C9_M7         Q9 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C9_M1         CONV_FLASH_C9_ND- N117007 CONV_FLASH_C9_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C9_M2         CONV_FLASH_C9_ND+ CONV_N117578 CONV_FLASH_C9_NDBIAS
+  0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C9_M3         CONV_FLASH_C9_ND- CONV_FLASH_C9_ND- N116990 N116990
+  CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_DECO_U31_M5         CONV_FLASH_DECO_ND2SB1 Q2 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U31_M6         CONV_FLASH_DECO_ND2SB1 Q2 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U16_M5         CONV_FLASH_DECO_N565094 Q16 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U16_M6         CONV_FLASH_DECO_N565094 Q16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U91_M5         CONV_FLASH_DECO_NDLSB16
+  CONV_FLASH_DECO_N578578 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U91_M6         CONV_FLASH_DECO_NDLSB16
+  CONV_FLASH_DECO_N578578 CONV_FLASH_DECO_U91_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U91_M2         CONV_FLASH_DECO_U91_ND2 Q31 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U91_M4         CONV_FLASH_DECO_NDLSB16 Q31 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U65_M5         CONV_FLASH_DECO_N568485
+  CONV_FLASH_DECO_N941987 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U65_M6         CONV_FLASH_DECO_N568485
+  CONV_FLASH_DECO_N941987 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U2_M5         CONV_FLASH_DECO_N259339 CONV_FLASH_D-MSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U2_M6         CONV_FLASH_DECO_N259339 CONV_FLASH_D-MSB 0 0
+  CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U96_M5         CONV_FLASH_DECO_NDLSB11
+  CONV_FLASH_DECO_N578514 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U96_M6         CONV_FLASH_DECO_NDLSB11
+  CONV_FLASH_DECO_N578514 CONV_FLASH_DECO_U96_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U96_M2         CONV_FLASH_DECO_U96_ND2 Q21 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U96_M4         CONV_FLASH_DECO_NDLSB11 Q21 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U109_M5         CONV_FLASH_DECO_N573020 Q48 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U109_M6         CONV_FLASH_DECO_N573020 Q48 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U57_M5         CONV_FLASH_DECO_ND2SB12
+  CONV_FLASH_DECO_N567821 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U57_M6         CONV_FLASH_DECO_ND2SB12
+  CONV_FLASH_DECO_N567821 CONV_FLASH_DECO_U57_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U57_M2         CONV_FLASH_DECO_U57_ND2 Q46 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U57_M4         CONV_FLASH_DECO_ND2SB12 Q46 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U28_M5         CONV_FLASH_DECO_ND3SB6 CONV_FLASH_DECO_N565120
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U28_M6         CONV_FLASH_DECO_ND3SB6 CONV_FLASH_DECO_N565120
+  CONV_FLASH_DECO_U28_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U28_M2         CONV_FLASH_DECO_U28_ND2 Q44 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U28_M4         CONV_FLASH_DECO_ND3SB6 Q44 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U139_M5         CONV_FLASH_DECO_NDX4LSB X4 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U139_M6         CONV_FLASH_DECO_NDX4LSB X4 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U74_M5         CONV_FLASH_DECO_N578674 Q12 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U74_M6         CONV_FLASH_DECO_N578674 Q12 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U43_M5         CONV_FLASH_DECO_N567821 Q44 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U43_M6         CONV_FLASH_DECO_N567821 Q44 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U80_M5         CONV_FLASH_DECO_N578524 Q22 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U80_M6         CONV_FLASH_DECO_N578524 Q22 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U14_M5         CONV_FLASH_DECO_ND3SB1 Q4 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U14_M6         CONV_FLASH_DECO_ND3SB1 Q4 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U136_M5         CONV_FLASH_DECO_NDX1LSB X1 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U136_M6         CONV_FLASH_DECO_NDX1LSB X1 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U124_M5         CONV_FLASH_DECO_NDLSB24
+  CONV_FLASH_DECO_N572160 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U124_M6         CONV_FLASH_DECO_NDLSB24
+  CONV_FLASH_DECO_N572160 CONV_FLASH_DECO_U124_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U124_M2         CONV_FLASH_DECO_U124_ND2 Q47 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U124_M4         CONV_FLASH_DECO_NDLSB24 Q47 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U116_M5         CONV_FLASH_DECO_N573096 Q62 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U116_M6         CONV_FLASH_DECO_N573096 Q62 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U69_M5         CONV_FLASH_DECO_N578608 Q2 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U69_M6         CONV_FLASH_DECO_N578608 Q2 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U86_M5         CONV_FLASH_DECO_NDLSB4 CONV_FLASH_DECO_N578636
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U86_M6         CONV_FLASH_DECO_NDLSB4 CONV_FLASH_DECO_N578636
+  CONV_FLASH_DECO_U86_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U86_M2         CONV_FLASH_DECO_U86_ND2 Q7 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U86_M4         CONV_FLASH_DECO_NDLSB4 Q7 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U26_M5         CONV_FLASH_DECO_ND3SB4 CONV_FLASH_DECO_N565104
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U26_M6         CONV_FLASH_DECO_ND3SB4 CONV_FLASH_DECO_N565104
+  CONV_FLASH_DECO_U26_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U26_M2         CONV_FLASH_DECO_U26_ND2 Q28 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U26_M4         CONV_FLASH_DECO_ND3SB4 Q28 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U103_M5         CONV_FLASH_DECO_N572104 Q36 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U103_M6         CONV_FLASH_DECO_N572104 Q36 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U37_M5         CONV_FLASH_DECO_N568555 Q24 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U37_M6         CONV_FLASH_DECO_N568555 Q24 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U61_M5         CONV_FLASH_DECO_ND2SB16
+  CONV_FLASH_DECO_N567861 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U61_M6         CONV_FLASH_DECO_ND2SB16
+  CONV_FLASH_DECO_N567861 CONV_FLASH_DECO_U61_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U61_M2         CONV_FLASH_DECO_U61_ND2 Q62 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U61_M4         CONV_FLASH_DECO_ND2SB16 Q62 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U119_M5         CONV_FLASH_DECO_NDLSB19
+  CONV_FLASH_DECO_N572104 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U119_M6         CONV_FLASH_DECO_NDLSB19
+  CONV_FLASH_DECO_N572104 CONV_FLASH_DECO_U119_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U119_M2         CONV_FLASH_DECO_U119_ND2 Q37 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U119_M4         CONV_FLASH_DECO_NDLSB19 Q37 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U48_M5         CONV_FLASH_DECO_ND2SB3 CONV_FLASH_DECO_N568511
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U48_M6         CONV_FLASH_DECO_ND2SB3 CONV_FLASH_DECO_N568511
+  CONV_FLASH_DECO_U48_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U48_M2         CONV_FLASH_DECO_U48_ND2 Q10 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U48_M4         CONV_FLASH_DECO_ND2SB3 Q10 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M16         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB12 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M5         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB16 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M11         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB9 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M9         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB14 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M1         CONV_FLASH_DECO_N941987 CONV_FLASH_DECO_ND2SB9
+  CONV_FLASH_DECO_U64_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M6         CONV_FLASH_DECO_U64_ND3
+  CONV_FLASH_DECO_ND2SB11 CONV_FLASH_DECO_U64_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M7         CONV_FLASH_DECO_U64_ND4
+  CONV_FLASH_DECO_ND2SB12 CONV_FLASH_DECO_U64_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M12         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB13 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M2         CONV_FLASH_DECO_U64_ND2
+  CONV_FLASH_DECO_ND2SB10 CONV_FLASH_DECO_U64_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M13         CONV_FLASH_DECO_U64_ND6
+  CONV_FLASH_DECO_ND2SB14 CONV_FLASH_DECO_U64_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M10         CONV_FLASH_DECO_U64_ND5
+  CONV_FLASH_DECO_ND2SB13 CONV_FLASH_DECO_U64_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M3         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB10 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M14         CONV_FLASH_DECO_U64_ND7
+  CONV_FLASH_DECO_ND2SB15 CONV_FLASH_DECO_U64_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U64_M8         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB15 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M4         CONV_FLASH_DECO_N941987
+  CONV_FLASH_DECO_ND2SB11 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U64_M15         CONV_FLASH_DECO_U64_ND8
+  CONV_FLASH_DECO_ND2SB16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U52_M5         CONV_FLASH_DECO_ND2SB7 CONV_FLASH_DECO_N568555
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U52_M6         CONV_FLASH_DECO_ND2SB7 CONV_FLASH_DECO_N568555
+  CONV_FLASH_DECO_U52_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U52_M2         CONV_FLASH_DECO_U52_ND2 Q26 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U52_M4         CONV_FLASH_DECO_ND2SB7 Q26 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U108_M5         CONV_FLASH_DECO_N572160 Q46 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U108_M6         CONV_FLASH_DECO_N572160 Q46 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U35_M5         CONV_FLASH_DECO_N568535 Q16 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U35_M6         CONV_FLASH_DECO_N568535 Q16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U24_M5         CONV_FLASH_DECO_ND3SB2 CONV_FLASH_DECO_N565082
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U24_M6         CONV_FLASH_DECO_ND3SB2 CONV_FLASH_DECO_N565082
+  CONV_FLASH_DECO_U24_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U24_M2         CONV_FLASH_DECO_U24_ND2 Q12 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U24_M4         CONV_FLASH_DECO_ND3SB2 Q12 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M16         X4 CONV_FLASH_DECO_NDLSB28 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M5         X4 CONV_FLASH_DECO_NDLSB32 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M11         X4 CONV_FLASH_DECO_NDLSB25 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M9         X4 CONV_FLASH_DECO_NDLSB30 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M1         X4 CONV_FLASH_DECO_NDLSB25
+  CONV_FLASH_DECO_U135_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M6         CONV_FLASH_DECO_U135_ND3
+  CONV_FLASH_DECO_NDLSB27 CONV_FLASH_DECO_U135_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M7         CONV_FLASH_DECO_U135_ND4
+  CONV_FLASH_DECO_NDLSB28 CONV_FLASH_DECO_U135_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M12         X4 CONV_FLASH_DECO_NDLSB29 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M2         CONV_FLASH_DECO_U135_ND2
+  CONV_FLASH_DECO_NDLSB26 CONV_FLASH_DECO_U135_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M13         CONV_FLASH_DECO_U135_ND6
+  CONV_FLASH_DECO_NDLSB30 CONV_FLASH_DECO_U135_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M10         CONV_FLASH_DECO_U135_ND5
+  CONV_FLASH_DECO_NDLSB29 CONV_FLASH_DECO_U135_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M3         X4 CONV_FLASH_DECO_NDLSB26 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M14         CONV_FLASH_DECO_U135_ND7
+  CONV_FLASH_DECO_NDLSB31 CONV_FLASH_DECO_U135_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U135_M8         X4 CONV_FLASH_DECO_NDLSB31 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M4         X4 CONV_FLASH_DECO_NDLSB27 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U135_M15         CONV_FLASH_DECO_U135_ND8
+  CONV_FLASH_DECO_NDLSB32 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U115_M5         CONV_FLASH_DECO_N573086 Q60 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U115_M6         CONV_FLASH_DECO_N573086 Q60 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U90_M5         CONV_FLASH_DECO_NDLSB8 CONV_FLASH_DECO_N578686
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U90_M6         CONV_FLASH_DECO_NDLSB8 CONV_FLASH_DECO_N578686
+  CONV_FLASH_DECO_U90_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U90_M2         CONV_FLASH_DECO_U90_ND2 Q15 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U90_M4         CONV_FLASH_DECO_NDLSB8 Q15 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U95_M5         CONV_FLASH_DECO_NDLSB12
+  CONV_FLASH_DECO_N578524 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U95_M6         CONV_FLASH_DECO_NDLSB12
+  CONV_FLASH_DECO_N578524 CONV_FLASH_DECO_U95_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U95_M2         CONV_FLASH_DECO_U95_ND2 Q23 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U95_M4         CONV_FLASH_DECO_NDLSB12 Q23 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U133_M5         CONV_FLASH_DECO_NDLSB25
+  CONV_FLASH_DECO_N573020 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U133_M6         CONV_FLASH_DECO_NDLSB25
+  CONV_FLASH_DECO_N573020 CONV_FLASH_DECO_U133_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U133_M2         CONV_FLASH_DECO_U133_ND2 Q49 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U133_M4         CONV_FLASH_DECO_NDLSB25 Q49 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U79_M5         CONV_FLASH_DECO_N578534 Q24 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U79_M6         CONV_FLASH_DECO_N578534 Q24 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U42_M5         CONV_FLASH_DECO_N567831 Q48 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U42_M6         CONV_FLASH_DECO_N567831 Q48 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U73_M5         CONV_FLASH_DECO_N578662 Q10 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U73_M6         CONV_FLASH_DECO_N578662 Q10 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U9_M5         CONV_FLASH_DECO_ND4SB3 CONV_FLASH_DECO_N259543
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U9_M6         CONV_FLASH_DECO_ND4SB3 CONV_FLASH_DECO_N259543
+  CONV_FLASH_DECO_U9_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U9_M2         CONV_FLASH_DECO_U9_ND2 Q40 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U9_M4         CONV_FLASH_DECO_ND4SB3 Q40 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U56_M5         CONV_FLASH_DECO_ND2SB11
+  CONV_FLASH_DECO_N567811 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U56_M6         CONV_FLASH_DECO_ND2SB11
+  CONV_FLASH_DECO_N567811 CONV_FLASH_DECO_U56_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U56_M2         CONV_FLASH_DECO_U56_ND2 Q42 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U56_M4         CONV_FLASH_DECO_ND2SB11 Q42 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U23_M5         CONV_FLASH_D-3SB CONV_FLASH_DECO_N565340
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U23_M6         CONV_FLASH_D-3SB CONV_FLASH_DECO_N565340 0 0
+  CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U123_M5         CONV_FLASH_DECO_NDLSB23
+  CONV_FLASH_DECO_N572144 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U123_M6         CONV_FLASH_DECO_NDLSB23
+  CONV_FLASH_DECO_N572144 CONV_FLASH_DECO_U123_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U123_M2         CONV_FLASH_DECO_U123_ND2 Q45 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U123_M4         CONV_FLASH_DECO_NDLSB23 Q45 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M16         CONV_FLASH_DECO_N567419
+  CONV_FLASH_DECO_ND2SB4 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M5         CONV_FLASH_DECO_N567419 CONV_FLASH_DECO_ND2SB8
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M11         CONV_FLASH_DECO_N567419
+  CONV_FLASH_DECO_ND2SB1 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M9         CONV_FLASH_DECO_N567419 CONV_FLASH_DECO_ND2SB6
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M1         CONV_FLASH_DECO_N567419 CONV_FLASH_DECO_ND2SB1
+  CONV_FLASH_DECO_U63_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M6         CONV_FLASH_DECO_U63_ND3 CONV_FLASH_DECO_ND2SB3
+  CONV_FLASH_DECO_U63_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M7         CONV_FLASH_DECO_U63_ND4 CONV_FLASH_DECO_ND2SB4
+  CONV_FLASH_DECO_U63_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M12         CONV_FLASH_DECO_N567419
+  CONV_FLASH_DECO_ND2SB5 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M2         CONV_FLASH_DECO_U63_ND2 CONV_FLASH_DECO_ND2SB2
+  CONV_FLASH_DECO_U63_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M13         CONV_FLASH_DECO_U63_ND6
+  CONV_FLASH_DECO_ND2SB6 CONV_FLASH_DECO_U63_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M10         CONV_FLASH_DECO_U63_ND5
+  CONV_FLASH_DECO_ND2SB5 CONV_FLASH_DECO_U63_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M3         CONV_FLASH_DECO_N567419 CONV_FLASH_DECO_ND2SB2
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M14         CONV_FLASH_DECO_U63_ND7
+  CONV_FLASH_DECO_ND2SB7 CONV_FLASH_DECO_U63_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U63_M8         CONV_FLASH_DECO_N567419 CONV_FLASH_DECO_ND2SB7
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M4         CONV_FLASH_DECO_N567419 CONV_FLASH_DECO_ND2SB3
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U63_M15         CONV_FLASH_DECO_U63_ND8
+  CONV_FLASH_DECO_ND2SB8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U21_M5         CONV_FLASH_DECO_N564924 Q56 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U21_M6         CONV_FLASH_DECO_N564924 Q56 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M16         X3 CONV_FLASH_DECO_NDLSB20 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M5         X3 CONV_FLASH_DECO_NDLSB24 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M11         X3 CONV_FLASH_DECO_NDLSB17 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M9         X3 CONV_FLASH_DECO_NDLSB22 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M1         X3 CONV_FLASH_DECO_NDLSB17
+  CONV_FLASH_DECO_U134_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M6         CONV_FLASH_DECO_U134_ND3
+  CONV_FLASH_DECO_NDLSB19 CONV_FLASH_DECO_U134_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M7         CONV_FLASH_DECO_U134_ND4
+  CONV_FLASH_DECO_NDLSB20 CONV_FLASH_DECO_U134_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M12         X3 CONV_FLASH_DECO_NDLSB21 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M2         CONV_FLASH_DECO_U134_ND2
+  CONV_FLASH_DECO_NDLSB18 CONV_FLASH_DECO_U134_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M13         CONV_FLASH_DECO_U134_ND6
+  CONV_FLASH_DECO_NDLSB22 CONV_FLASH_DECO_U134_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M10         CONV_FLASH_DECO_U134_ND5
+  CONV_FLASH_DECO_NDLSB21 CONV_FLASH_DECO_U134_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M3         X3 CONV_FLASH_DECO_NDLSB18 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M14         CONV_FLASH_DECO_U134_ND7
+  CONV_FLASH_DECO_NDLSB23 CONV_FLASH_DECO_U134_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U134_M8         X3 CONV_FLASH_DECO_NDLSB23 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M4         X3 CONV_FLASH_DECO_NDLSB19 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U134_M15         CONV_FLASH_DECO_U134_ND8
+  CONV_FLASH_DECO_NDLSB24 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U3_M5         CONV_FLASH_DECO_N259565 Q16 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U3_M6         CONV_FLASH_DECO_N259565 Q16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U114_M5         CONV_FLASH_DECO_N573076 Q58 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U114_M6         CONV_FLASH_DECO_N573076 Q58 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U6_M5         CONV_FLASH_D-5SB CONV_FLASH_DECO_ND5SB1 N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U6_M6         CONV_FLASH_D-5SB CONV_FLASH_DECO_ND5SB1
+  CONV_FLASH_DECO_U6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U6_M2         CONV_FLASH_DECO_U6_ND2 CONV_FLASH_DECO_ND5SB2 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U6_M4         CONV_FLASH_D-5SB CONV_FLASH_DECO_ND5SB2 N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U102_M5         CONV_FLASH_DECO_N572074 Q34 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U102_M6         CONV_FLASH_DECO_N572074 Q34 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U36_M5         CONV_FLASH_DECO_N568545 Q20 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U36_M6         CONV_FLASH_DECO_N568545 Q20 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U68_M5         CONV_FLASH_DECO_NDLSB1 Q1 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U68_M6         CONV_FLASH_DECO_NDLSB1 Q1 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U85_M5         CONV_FLASH_DECO_NDLSB3 CONV_FLASH_DECO_N578622
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U85_M6         CONV_FLASH_DECO_NDLSB3 CONV_FLASH_DECO_N578622
+  CONV_FLASH_DECO_U85_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U85_M2         CONV_FLASH_DECO_U85_ND2 Q5 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U85_M4         CONV_FLASH_DECO_NDLSB3 Q5 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U107_M5         CONV_FLASH_DECO_N572144 Q44 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U107_M6         CONV_FLASH_DECO_N572144 Q44 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U140_M7         CONV_FLASH_D-LSB CONV_FLASH_DECO_NDX1LSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U140_M8         CONV_FLASH_D-LSB CONV_FLASH_DECO_NDX2LSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U140_M12         CONV_FLASH_D-LSB CONV_FLASH_DECO_NDX4LSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U140_M9         CONV_FLASH_D-LSB CONV_FLASH_DECO_NDX3LSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U140_M1         CONV_FLASH_D-LSB CONV_FLASH_DECO_NDX1LSB
+  CONV_FLASH_DECO_U140_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U140_M10         CONV_FLASH_DECO_U140_ND3
+  CONV_FLASH_DECO_NDX3LSB CONV_FLASH_DECO_U140_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U140_M3         CONV_FLASH_DECO_U140_ND2
+  CONV_FLASH_DECO_NDX2LSB CONV_FLASH_DECO_U140_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U140_M11         CONV_FLASH_DECO_U140_ND4
+  CONV_FLASH_DECO_NDX4LSB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U78_M5         CONV_FLASH_DECO_N578552 Q26 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U78_M6         CONV_FLASH_DECO_N578552 Q26 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U60_M5         CONV_FLASH_DECO_ND2SB15
+  CONV_FLASH_DECO_N567851 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U60_M6         CONV_FLASH_DECO_ND2SB15
+  CONV_FLASH_DECO_N567851 CONV_FLASH_DECO_U60_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U60_M2         CONV_FLASH_DECO_U60_ND2 Q58 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U60_M4         CONV_FLASH_DECO_ND2SB15 Q58 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U120_M5         CONV_FLASH_DECO_NDLSB20
+  CONV_FLASH_DECO_N793529 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U120_M6         CONV_FLASH_DECO_NDLSB20
+  CONV_FLASH_DECO_N793529 CONV_FLASH_DECO_U120_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U120_M2         CONV_FLASH_DECO_U120_ND2 Q39 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U120_M4         CONV_FLASH_DECO_NDLSB20 Q39 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U19_M5         CONV_FLASH_DECO_N565120 Q40 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U19_M6         CONV_FLASH_DECO_N565120 Q40 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U41_M5         CONV_FLASH_DECO_N567841 Q52 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U41_M6         CONV_FLASH_DECO_N567841 Q52 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U118_M5         CONV_FLASH_DECO_NDLSB18
+  CONV_FLASH_DECO_N572074 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U118_M6         CONV_FLASH_DECO_NDLSB18
+  CONV_FLASH_DECO_N572074 CONV_FLASH_DECO_U118_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U118_M2         CONV_FLASH_DECO_U118_ND2 Q35 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U118_M4         CONV_FLASH_DECO_NDLSB18 Q35 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U132_M5         CONV_FLASH_DECO_NDLSB26
+  CONV_FLASH_DECO_N573036 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U132_M6         CONV_FLASH_DECO_NDLSB26
+  CONV_FLASH_DECO_N573036 CONV_FLASH_DECO_U132_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U132_M2         CONV_FLASH_DECO_U132_ND2 Q51 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U132_M4         CONV_FLASH_DECO_NDLSB26 Q51 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U34_M5         CONV_FLASH_DECO_N568523 Q12 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U34_M6         CONV_FLASH_DECO_N568523 Q12 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U137_M5         CONV_FLASH_DECO_NDX2LSB X2 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U137_M6         CONV_FLASH_DECO_NDX2LSB X2 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U94_M5         CONV_FLASH_DECO_NDLSB13
+  CONV_FLASH_DECO_N578534 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U94_M6         CONV_FLASH_DECO_NDLSB13
+  CONV_FLASH_DECO_N578534 CONV_FLASH_DECO_U94_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U94_M2         CONV_FLASH_DECO_U94_ND2 Q25 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U94_M4         CONV_FLASH_DECO_NDLSB13 Q25 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U51_M5         CONV_FLASH_DECO_ND2SB6 CONV_FLASH_DECO_N568545
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U51_M6         CONV_FLASH_DECO_ND2SB6 CONV_FLASH_DECO_N568545
+  CONV_FLASH_DECO_U51_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U51_M2         CONV_FLASH_DECO_U51_ND2 Q22 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U51_M4         CONV_FLASH_DECO_ND2SB6 Q22 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U89_M5         CONV_FLASH_DECO_NDLSB7 CONV_FLASH_DECO_N578674
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U89_M6         CONV_FLASH_DECO_NDLSB7 CONV_FLASH_DECO_N578674
+  CONV_FLASH_DECO_U89_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U89_M2         CONV_FLASH_DECO_U89_ND2 Q13 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U89_M4         CONV_FLASH_DECO_NDLSB7 Q13 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U47_M5         CONV_FLASH_DECO_ND2SB2 CONV_FLASH_DECO_N568499
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U47_M6         CONV_FLASH_DECO_ND2SB2 CONV_FLASH_DECO_N568499
+  CONV_FLASH_DECO_U47_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U47_M2         CONV_FLASH_DECO_U47_ND2 Q6 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U47_M4         CONV_FLASH_DECO_ND2SB2 Q6 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U72_M5         CONV_FLASH_DECO_N578650 Q8 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U72_M6         CONV_FLASH_DECO_N578650 Q8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U17_M5         CONV_FLASH_DECO_N565104 Q24 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U17_M6         CONV_FLASH_DECO_N565104 Q24 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U113_M5         CONV_FLASH_DECO_N573066 Q56 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U113_M6         CONV_FLASH_DECO_N573066 Q56 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M16         X2 CONV_FLASH_DECO_NDLSB12 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M5         X2 CONV_FLASH_DECO_NDLSB16 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M11         X2 CONV_FLASH_DECO_NDLSB9 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M9         X2 CONV_FLASH_DECO_NDLSB14 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M1         X2 CONV_FLASH_DECO_NDLSB9
+  CONV_FLASH_DECO_U100_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M6         CONV_FLASH_DECO_U100_ND3
+  CONV_FLASH_DECO_NDLSB11 CONV_FLASH_DECO_U100_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M7         CONV_FLASH_DECO_U100_ND4
+  CONV_FLASH_DECO_NDLSB12 CONV_FLASH_DECO_U100_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M12         X2 CONV_FLASH_DECO_NDLSB13 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M2         CONV_FLASH_DECO_U100_ND2
+  CONV_FLASH_DECO_NDLSB10 CONV_FLASH_DECO_U100_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M13         CONV_FLASH_DECO_U100_ND6
+  CONV_FLASH_DECO_NDLSB14 CONV_FLASH_DECO_U100_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M10         CONV_FLASH_DECO_U100_ND5
+  CONV_FLASH_DECO_NDLSB13 CONV_FLASH_DECO_U100_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M3         X2 CONV_FLASH_DECO_NDLSB10 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M14         CONV_FLASH_DECO_U100_ND7
+  CONV_FLASH_DECO_NDLSB15 CONV_FLASH_DECO_U100_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U100_M8         X2 CONV_FLASH_DECO_NDLSB15 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M4         X2 CONV_FLASH_DECO_NDLSB11 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U100_M15         CONV_FLASH_DECO_U100_ND8
+  CONV_FLASH_DECO_NDLSB16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U55_M5         CONV_FLASH_DECO_ND2SB10
+  CONV_FLASH_DECO_N567801 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U55_M6         CONV_FLASH_DECO_ND2SB10
+  CONV_FLASH_DECO_N567801 CONV_FLASH_DECO_U55_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U55_M2         CONV_FLASH_DECO_U55_ND2 Q38 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U55_M4         CONV_FLASH_DECO_ND2SB10 Q38 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U29_M5         CONV_FLASH_DECO_ND3SB7 CONV_FLASH_DECO_N565130
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U29_M6         CONV_FLASH_DECO_ND3SB7 CONV_FLASH_DECO_N565130
+  CONV_FLASH_DECO_U29_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U29_M2         CONV_FLASH_DECO_U29_ND2 Q52 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U29_M4         CONV_FLASH_DECO_ND3SB7 Q52 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U127_M5         CONV_FLASH_DECO_NDLSB30
+  CONV_FLASH_DECO_N573076 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U127_M6         CONV_FLASH_DECO_NDLSB30
+  CONV_FLASH_DECO_N573076 CONV_FLASH_DECO_U127_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U127_M2         CONV_FLASH_DECO_U127_ND2 Q59 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U127_M4         CONV_FLASH_DECO_NDLSB30 Q59 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U122_M5         CONV_FLASH_DECO_NDLSB22
+  CONV_FLASH_DECO_N572134 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U122_M6         CONV_FLASH_DECO_NDLSB22
+  CONV_FLASH_DECO_N572134 CONV_FLASH_DECO_U122_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U122_M2         CONV_FLASH_DECO_U122_ND2 Q43 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U122_M4         CONV_FLASH_DECO_NDLSB22 Q43 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U106_M5         CONV_FLASH_DECO_N572134 Q42 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U106_M6         CONV_FLASH_DECO_N572134 Q42 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U77_M5         CONV_FLASH_DECO_N578562 Q28 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U77_M6         CONV_FLASH_DECO_N578562 Q28 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U15_M5         CONV_FLASH_DECO_N565082 Q8 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U15_M6         CONV_FLASH_DECO_N565082 Q8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U10_M5         CONV_FLASH_DECO_ND4SB4 CONV_FLASH_DECO_N259605
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U10_M6         CONV_FLASH_DECO_ND4SB4 CONV_FLASH_DECO_N259605
+  CONV_FLASH_DECO_U10_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U10_M2         CONV_FLASH_DECO_U10_ND2 Q56 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U10_M4         CONV_FLASH_DECO_ND4SB4 Q56 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U40_M5         CONV_FLASH_DECO_N567851 Q56 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U40_M6         CONV_FLASH_DECO_N567851 Q56 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U131_M5         CONV_FLASH_DECO_NDLSB27
+  CONV_FLASH_DECO_N573046 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U131_M6         CONV_FLASH_DECO_NDLSB27
+  CONV_FLASH_DECO_N573046 CONV_FLASH_DECO_U131_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U131_M2         CONV_FLASH_DECO_U131_ND2 Q53 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U131_M4         CONV_FLASH_DECO_NDLSB27 Q53 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U101_M5         CONV_FLASH_DECO_N572064 CONV_FLASH_D-MSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U101_M6         CONV_FLASH_DECO_N572064 CONV_FLASH_D-MSB 0 0
+  CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U27_M5         CONV_FLASH_DECO_ND3SB5 CONV_FLASH_DECO_N564920
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U27_M6         CONV_FLASH_DECO_ND3SB5 CONV_FLASH_DECO_N564920
+  CONV_FLASH_DECO_U27_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U27_M2         CONV_FLASH_DECO_U27_ND2 Q36 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U27_M4         CONV_FLASH_DECO_ND3SB5 Q36 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U84_M5         CONV_FLASH_DECO_NDLSB2 CONV_FLASH_DECO_N578608
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U84_M6         CONV_FLASH_DECO_NDLSB2 CONV_FLASH_DECO_N578608
+  CONV_FLASH_DECO_U84_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U84_M2         CONV_FLASH_DECO_U84_ND2 Q3 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U84_M4         CONV_FLASH_DECO_NDLSB2 Q3 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U59_M5         CONV_FLASH_DECO_ND2SB14
+  CONV_FLASH_DECO_N567841 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U59_M6         CONV_FLASH_DECO_ND2SB14
+  CONV_FLASH_DECO_N567841 CONV_FLASH_DECO_U59_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U59_M2         CONV_FLASH_DECO_U59_ND2 Q54 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U59_M4         CONV_FLASH_DECO_ND2SB14 Q54 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M16         CONV_FLASH_DECO_N565498
+  CONV_FLASH_DECO_ND3SB4 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M5         CONV_FLASH_DECO_N565498 CONV_FLASH_DECO_ND3SB8
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M11         CONV_FLASH_DECO_N565498
+  CONV_FLASH_DECO_ND3SB1 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M9         CONV_FLASH_DECO_N565498 CONV_FLASH_DECO_ND3SB6
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M1         CONV_FLASH_DECO_N565498 CONV_FLASH_DECO_ND3SB1
+  CONV_FLASH_DECO_U13_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M6         CONV_FLASH_DECO_U13_ND3 CONV_FLASH_DECO_ND3SB3
+  CONV_FLASH_DECO_U13_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M7         CONV_FLASH_DECO_U13_ND4 CONV_FLASH_DECO_ND3SB4
+  CONV_FLASH_DECO_U13_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M12         CONV_FLASH_DECO_N565498
+  CONV_FLASH_DECO_ND3SB5 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M2         CONV_FLASH_DECO_U13_ND2 CONV_FLASH_DECO_ND3SB2
+  CONV_FLASH_DECO_U13_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M13         CONV_FLASH_DECO_U13_ND6
+  CONV_FLASH_DECO_ND3SB6 CONV_FLASH_DECO_U13_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M10         CONV_FLASH_DECO_U13_ND5
+  CONV_FLASH_DECO_ND3SB5 CONV_FLASH_DECO_U13_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M3         CONV_FLASH_DECO_N565498 CONV_FLASH_DECO_ND3SB2
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M14         CONV_FLASH_DECO_U13_ND7
+  CONV_FLASH_DECO_ND3SB7 CONV_FLASH_DECO_U13_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U13_M8         CONV_FLASH_DECO_N565498 CONV_FLASH_DECO_ND3SB7
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M4         CONV_FLASH_DECO_N565498 CONV_FLASH_DECO_ND3SB3
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U13_M15         CONV_FLASH_DECO_U13_ND8
+  CONV_FLASH_DECO_ND3SB8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U112_M5         CONV_FLASH_DECO_N573056 Q54 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U112_M6         CONV_FLASH_DECO_N573056 Q54 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U93_M5         CONV_FLASH_DECO_NDLSB14
+  CONV_FLASH_DECO_N578552 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U93_M6         CONV_FLASH_DECO_NDLSB14
+  CONV_FLASH_DECO_N578552 CONV_FLASH_DECO_U93_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U93_M2         CONV_FLASH_DECO_U93_ND2 Q27 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U93_M4         CONV_FLASH_DECO_NDLSB14 Q27 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M16         X1 CONV_FLASH_DECO_NDLSB4 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M5         X1 CONV_FLASH_DECO_NDLSB8 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M11         X1 CONV_FLASH_DECO_NDLSB1 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M9         X1 CONV_FLASH_DECO_NDLSB6 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M1         X1 CONV_FLASH_DECO_NDLSB1
+  CONV_FLASH_DECO_U99_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M6         CONV_FLASH_DECO_U99_ND3 CONV_FLASH_DECO_NDLSB3
+  CONV_FLASH_DECO_U99_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M7         CONV_FLASH_DECO_U99_ND4 CONV_FLASH_DECO_NDLSB4
+  CONV_FLASH_DECO_U99_ND5 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M12         X1 CONV_FLASH_DECO_NDLSB5 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M2         CONV_FLASH_DECO_U99_ND2 CONV_FLASH_DECO_NDLSB2
+  CONV_FLASH_DECO_U99_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M13         CONV_FLASH_DECO_U99_ND6
+  CONV_FLASH_DECO_NDLSB6 CONV_FLASH_DECO_U99_ND7 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M10         CONV_FLASH_DECO_U99_ND5
+  CONV_FLASH_DECO_NDLSB5 CONV_FLASH_DECO_U99_ND6 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M3         X1 CONV_FLASH_DECO_NDLSB2 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M14         CONV_FLASH_DECO_U99_ND7
+  CONV_FLASH_DECO_NDLSB7 CONV_FLASH_DECO_U99_ND8 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U99_M8         X1 CONV_FLASH_DECO_NDLSB7 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M4         X1 CONV_FLASH_DECO_NDLSB3 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U99_M15         CONV_FLASH_DECO_U99_ND8
+  CONV_FLASH_DECO_NDLSB8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U117_M5         CONV_FLASH_DECO_NDLSB17
+  CONV_FLASH_DECO_N572064 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U117_M6         CONV_FLASH_DECO_NDLSB17
+  CONV_FLASH_DECO_N572064 CONV_FLASH_DECO_U117_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U117_M2         CONV_FLASH_DECO_U117_ND2 Q33 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U117_M4         CONV_FLASH_DECO_NDLSB17 Q33 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U33_M5         CONV_FLASH_DECO_N568511 Q8 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U33_M6         CONV_FLASH_DECO_N568511 Q8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U98_M5         CONV_FLASH_DECO_NDLSB9 CONV_FLASH_DECO_N578480
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U98_M6         CONV_FLASH_DECO_NDLSB9 CONV_FLASH_DECO_N578480
+  CONV_FLASH_DECO_U98_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U98_M2         CONV_FLASH_DECO_U98_ND2 Q17 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U98_M4         CONV_FLASH_DECO_NDLSB9 Q17 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U4_M5         CONV_FLASH_DECO_N259543 CONV_FLASH_D-MSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U4_M6         CONV_FLASH_DECO_N259543 CONV_FLASH_D-MSB 0 0
+  CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U46_M5         CONV_FLASH_DECO_N569141 CONV_FLASH_D-MSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U46_M6         CONV_FLASH_DECO_N569141 CONV_FLASH_D-MSB 0 0
+  CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U7_M5         CONV_FLASH_DECO_ND5SB2 CONV_FLASH_DECO_N259339
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U7_M6         CONV_FLASH_DECO_ND5SB2 CONV_FLASH_DECO_N259339
+  CONV_FLASH_DECO_U7_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U7_M2         CONV_FLASH_DECO_U7_ND2 Q48 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U7_M4         CONV_FLASH_DECO_ND5SB2 Q48 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U71_M5         CONV_FLASH_DECO_N578636 Q6 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U71_M6         CONV_FLASH_DECO_N578636 Q6 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U88_M5         CONV_FLASH_DECO_NDLSB6 CONV_FLASH_DECO_N578662
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U88_M6         CONV_FLASH_DECO_NDLSB6 CONV_FLASH_DECO_N578662
+  CONV_FLASH_DECO_U88_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U88_M2         CONV_FLASH_DECO_U88_ND2 Q11 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U88_M4         CONV_FLASH_DECO_NDLSB6 Q11 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U25_M5         CONV_FLASH_DECO_ND3SB3 CONV_FLASH_DECO_N565094
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U25_M6         CONV_FLASH_DECO_ND3SB3 CONV_FLASH_DECO_N565094
+  CONV_FLASH_DECO_U25_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U25_M2         CONV_FLASH_DECO_U25_ND2 Q20 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U25_M4         CONV_FLASH_DECO_ND3SB3 Q20 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U50_M5         CONV_FLASH_DECO_ND2SB5 CONV_FLASH_DECO_N568535
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U50_M6         CONV_FLASH_DECO_ND2SB5 CONV_FLASH_DECO_N568535
+  CONV_FLASH_DECO_U50_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U50_M2         CONV_FLASH_DECO_U50_ND2 Q18 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U50_M4         CONV_FLASH_DECO_ND2SB5 Q18 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U76_M5         CONV_FLASH_DECO_N578578 Q30 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U76_M6         CONV_FLASH_DECO_N578578 Q30 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U126_M5         CONV_FLASH_DECO_NDLSB31
+  CONV_FLASH_DECO_N573086 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U126_M6         CONV_FLASH_DECO_NDLSB31
+  CONV_FLASH_DECO_N573086 CONV_FLASH_DECO_U126_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U126_M2         CONV_FLASH_DECO_U126_ND2 Q61 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U126_M4         CONV_FLASH_DECO_NDLSB31 Q61 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U1_M5         CONV_FLASH_DECO_ND5SB1 Q16 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U1_M6         CONV_FLASH_DECO_ND5SB1 Q16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U105_M5         CONV_FLASH_DECO_N572124 Q40 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U105_M6         CONV_FLASH_DECO_N572124 Q40 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U83_M5         CONV_FLASH_DECO_N578480 Q16 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U83_M6         CONV_FLASH_DECO_N578480 Q16 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U54_M5         CONV_FLASH_DECO_ND2SB9 CONV_FLASH_DECO_N569141
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U54_M6         CONV_FLASH_DECO_ND2SB9 CONV_FLASH_DECO_N569141
+  CONV_FLASH_DECO_U54_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U54_M2         CONV_FLASH_DECO_U54_ND2 Q34 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U54_M4         CONV_FLASH_DECO_ND2SB9 Q34 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U12_M7         CONV_FLASH_D-4SB CONV_FLASH_DECO_ND4SB1
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U12_M8         CONV_FLASH_D-4SB CONV_FLASH_DECO_ND4SB2
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U12_M12         CONV_FLASH_D-4SB CONV_FLASH_DECO_ND4SB4
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U12_M9         CONV_FLASH_D-4SB CONV_FLASH_DECO_ND4SB3
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U12_M1         CONV_FLASH_D-4SB CONV_FLASH_DECO_ND4SB1
+  CONV_FLASH_DECO_U12_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U12_M10         CONV_FLASH_DECO_U12_ND3
+  CONV_FLASH_DECO_ND4SB3 CONV_FLASH_DECO_U12_ND4 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U12_M3         CONV_FLASH_DECO_U12_ND2 CONV_FLASH_DECO_ND4SB2
+  CONV_FLASH_DECO_U12_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U12_M11         CONV_FLASH_DECO_U12_ND4
+  CONV_FLASH_DECO_ND4SB4 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U138_M5         CONV_FLASH_DECO_NDX3LSB X3 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U138_M6         CONV_FLASH_DECO_NDX3LSB X3 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U121_M5         CONV_FLASH_DECO_NDLSB21
+  CONV_FLASH_DECO_N572124 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U121_M6         CONV_FLASH_DECO_NDLSB21
+  CONV_FLASH_DECO_N572124 CONV_FLASH_DECO_U121_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U121_M2         CONV_FLASH_DECO_U121_ND2 Q41 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U121_M4         CONV_FLASH_DECO_NDLSB21 Q41 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U111_M5         CONV_FLASH_DECO_N573046 Q52 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U111_M6         CONV_FLASH_DECO_N573046 Q52 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U130_M5         CONV_FLASH_DECO_NDLSB28
+  CONV_FLASH_DECO_N573056 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U130_M6         CONV_FLASH_DECO_NDLSB28
+  CONV_FLASH_DECO_N573056 CONV_FLASH_DECO_U130_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U130_M2         CONV_FLASH_DECO_U130_ND2 Q55 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U130_M4         CONV_FLASH_DECO_NDLSB28 Q55 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U39_M5         CONV_FLASH_DECO_N567861 Q60 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U39_M6         CONV_FLASH_DECO_N567861 Q60 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U30_M5         CONV_FLASH_DECO_ND3SB8 CONV_FLASH_DECO_N564924
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U30_M6         CONV_FLASH_DECO_ND3SB8 CONV_FLASH_DECO_N564924
+  CONV_FLASH_DECO_U30_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U30_M2         CONV_FLASH_DECO_U30_ND2 Q60 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U30_M4         CONV_FLASH_DECO_ND3SB8 Q60 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U45_M5         CONV_FLASH_DECO_N567801 Q36 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U45_M6         CONV_FLASH_DECO_N567801 Q36 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U22_M5         CONV_FLASH_DECO_N565340
+  CONV_FLASH_DECO_N565498 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U22_M6         CONV_FLASH_DECO_N565340
+  CONV_FLASH_DECO_N565498 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U92_M5         CONV_FLASH_DECO_NDLSB15
+  CONV_FLASH_DECO_N578562 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U92_M6         CONV_FLASH_DECO_NDLSB15
+  CONV_FLASH_DECO_N578562 CONV_FLASH_DECO_U92_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U92_M2         CONV_FLASH_DECO_U92_ND2 Q29 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U92_M4         CONV_FLASH_DECO_NDLSB15 Q29 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U58_M5         CONV_FLASH_DECO_ND2SB13
+  CONV_FLASH_DECO_N567831 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U58_M6         CONV_FLASH_DECO_ND2SB13
+  CONV_FLASH_DECO_N567831 CONV_FLASH_DECO_U58_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U58_M2         CONV_FLASH_DECO_U58_ND2 Q50 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U58_M4         CONV_FLASH_DECO_ND2SB13 Q50 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U97_M5         CONV_FLASH_DECO_NDLSB10
+  CONV_FLASH_DECO_N578504 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U97_M6         CONV_FLASH_DECO_NDLSB10
+  CONV_FLASH_DECO_N578504 CONV_FLASH_DECO_U97_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U97_M2         CONV_FLASH_DECO_U97_ND2 Q19 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U97_M4         CONV_FLASH_DECO_NDLSB10 Q19 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U82_M5         CONV_FLASH_DECO_N578504 Q18 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U82_M6         CONV_FLASH_DECO_N578504 Q18 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U20_M5         CONV_FLASH_DECO_N565130 Q48 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U20_M6         CONV_FLASH_DECO_N565130 Q48 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U32_M5         CONV_FLASH_DECO_N568499 Q4 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U32_M6         CONV_FLASH_DECO_N568499 Q4 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U75_M5         CONV_FLASH_DECO_N578686 Q14 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U75_M6         CONV_FLASH_DECO_N578686 Q14 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U70_M5         CONV_FLASH_DECO_N578622 Q4 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U70_M6         CONV_FLASH_DECO_N578622 Q4 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U87_M5         CONV_FLASH_DECO_NDLSB5 CONV_FLASH_DECO_N578650
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U87_M6         CONV_FLASH_DECO_NDLSB5 CONV_FLASH_DECO_N578650
+  CONV_FLASH_DECO_U87_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U87_M2         CONV_FLASH_DECO_U87_ND2 Q9 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U87_M4         CONV_FLASH_DECO_NDLSB5 Q9 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U110_M5         CONV_FLASH_DECO_N573036 Q50 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U110_M6         CONV_FLASH_DECO_N573036 Q50 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U125_M5         CONV_FLASH_DECO_NDLSB32
+  CONV_FLASH_DECO_N573096 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U125_M6         CONV_FLASH_DECO_NDLSB32
+  CONV_FLASH_DECO_N573096 CONV_FLASH_DECO_U125_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U125_M2         CONV_FLASH_DECO_U125_ND2 Q63 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U125_M4         CONV_FLASH_DECO_NDLSB32 Q63 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U67_M5         CONV_FLASH_DECO_N567401
+  CONV_FLASH_DECO_N567419 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U67_M6         CONV_FLASH_DECO_N567401
+  CONV_FLASH_DECO_N567419 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U11_M5         CONV_FLASH_DECO_ND4SB1 Q8 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U11_M6         CONV_FLASH_DECO_ND4SB1 Q8 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U49_M5         CONV_FLASH_DECO_ND2SB4 CONV_FLASH_DECO_N568523
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U49_M6         CONV_FLASH_DECO_ND2SB4 CONV_FLASH_DECO_N568523
+  CONV_FLASH_DECO_U49_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U49_M2         CONV_FLASH_DECO_U49_ND2 Q14 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U49_M4         CONV_FLASH_DECO_ND2SB4 Q14 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U104_M5         CONV_FLASH_DECO_N793529 Q38 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U104_M6         CONV_FLASH_DECO_N793529 Q38 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U18_M5         CONV_FLASH_DECO_N564920 CONV_FLASH_D-MSB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U18_M6         CONV_FLASH_DECO_N564920 CONV_FLASH_D-MSB 0 0
+  CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U129_M5         CONV_FLASH_DECO_NDLSB29
+  CONV_FLASH_DECO_N573066 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U129_M6         CONV_FLASH_DECO_NDLSB29
+  CONV_FLASH_DECO_N573066 CONV_FLASH_DECO_U129_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U129_M2         CONV_FLASH_DECO_U129_ND2 Q57 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U129_M4         CONV_FLASH_DECO_NDLSB29 Q57 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U44_M5         CONV_FLASH_DECO_N567811 Q40 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U44_M6         CONV_FLASH_DECO_N567811 Q40 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U38_M5         CONV_FLASH_DECO_N568565 Q28 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U38_M6         CONV_FLASH_DECO_N568565 Q28 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U53_M5         CONV_FLASH_DECO_ND2SB8 CONV_FLASH_DECO_N568565
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U53_M6         CONV_FLASH_DECO_ND2SB8 CONV_FLASH_DECO_N568565
+  CONV_FLASH_DECO_U53_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U53_M2         CONV_FLASH_DECO_U53_ND2 Q30 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U53_M4         CONV_FLASH_DECO_ND2SB8 Q30 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U8_M5         CONV_FLASH_DECO_ND4SB2 CONV_FLASH_DECO_N259565
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U8_M6         CONV_FLASH_DECO_ND4SB2 CONV_FLASH_DECO_N259565
+  CONV_FLASH_DECO_U8_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U8_M2         CONV_FLASH_DECO_U8_ND2 Q24 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U8_M4         CONV_FLASH_DECO_ND4SB2 Q24 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U62_M5         CONV_FLASH_D-2SB CONV_FLASH_DECO_N568485
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U62_M6         CONV_FLASH_D-2SB CONV_FLASH_DECO_N568485
+  CONV_FLASH_DECO_U62_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U62_M2         CONV_FLASH_DECO_U62_ND2
+  CONV_FLASH_DECO_N567401 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U62_M4         CONV_FLASH_D-2SB CONV_FLASH_DECO_N567401
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U5_M5         CONV_FLASH_DECO_N259605 Q48 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U5_M6         CONV_FLASH_DECO_N259605 Q48 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_DECO_U81_M5         CONV_FLASH_DECO_N578514 Q20 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_DECO_U81_M6         CONV_FLASH_DECO_N578514 Q20 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_C24_M4         CONV_FLASH_C24_ND+ CONV_FLASH_C24_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C24_M5         CONV_FLASH_C24_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C24_M6         Q24 CONV_FLASH_C24_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C24_M7         Q24 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C24_M1         CONV_FLASH_C24_ND- N117007 CONV_FLASH_C24_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C24_M2         CONV_FLASH_C24_ND+ CONV_N117532
+  CONV_FLASH_C24_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C24_M3         CONV_FLASH_C24_ND- CONV_FLASH_C24_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_FFD2_NAND6_M5         CONV_FLASH_FFD2_N62152 CONV_FLASH_FFD2_Y
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND6_M6         CONV_FLASH_FFD2_N62152 CONV_FLASH_FFD2_Y
+  CONV_FLASH_FFD2_NAND6_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND6_M2         CONV_FLASH_FFD2_NAND6_ND2 CONV_FLASH_D-2SB 0
+  0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND6_M4         CONV_FLASH_FFD2_N62152 CONV_FLASH_D-2SB
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND1_M2         CONV_FLASH_FFD2_NAND1_ND2 N116976
+  CONV_FLASH_FFD2_NAND1_ND3 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND1_M3         CONV_FLASH_FFD2_Y CONV_FLASH_FFD2_X N116990
+  N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND1_M6         CONV_FLASH_FFD2_NAND1_ND3
+  CONV_FLASH_FFD2_N62152 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND1_M4         CONV_FLASH_FFD2_Y N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND1_M1         CONV_FLASH_FFD2_Y CONV_FLASH_FFD2_X
+  CONV_FLASH_FFD2_NAND1_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND1_M5         CONV_FLASH_FFD2_Y CONV_FLASH_FFD2_N62152
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND2_M5         CONV_FLASH_FFD2_N62128
+  CONV_FLASH_FFD2_N62152 N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND2_M6         CONV_FLASH_FFD2_N62128
+  CONV_FLASH_FFD2_N62152 CONV_FLASH_FFD2_NAND2_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND2_M2         CONV_FLASH_FFD2_NAND2_ND2 CONV_FLASH_FFD2_X
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND2_M4         CONV_FLASH_FFD2_N62128 CONV_FLASH_FFD2_X
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND3_M5         CONV_FLASH_FFD2_X CONV_FLASH_FFD2_N62128
+  N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND3_M6         CONV_FLASH_FFD2_X CONV_FLASH_FFD2_N62128
+  CONV_FLASH_FFD2_NAND3_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND3_M2         CONV_FLASH_FFD2_NAND3_ND2 N116976 0 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND3_M4         CONV_FLASH_FFD2_X N116976 N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND4_M5         2SB CONV_FLASH_FFD2_X N116990 N116990 CMOSP 
+  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND4_M6         2SB CONV_FLASH_FFD2_X
+  CONV_FLASH_FFD2_NAND4_ND2 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND4_M2         CONV_FLASH_FFD2_NAND4_ND2 N-2SB 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND4_M4         2SB N-2SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND5_M5         N-2SB 2SB N116990 N116990 CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_FFD2_NAND5_M6         N-2SB 2SB CONV_FLASH_FFD2_NAND5_ND2 0 CMOSN 
+  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND5_M2         CONV_FLASH_FFD2_NAND5_ND2 CONV_FLASH_FFD2_Y
+  0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_CONV_FLASH_FFD2_NAND5_M4         N-2SB CONV_FLASH_FFD2_Y N116990 N116990
+  CMOSP  
+ L=.18u  
+ W=.2u         
M_CONV_FLASH_C20_M4         CONV_FLASH_C20_ND+ CONV_FLASH_C20_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C20_M5         CONV_FLASH_C20_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C20_M6         Q20 CONV_FLASH_C20_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C20_M7         Q20 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C20_M1         CONV_FLASH_C20_ND- N117007 CONV_FLASH_C20_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C20_M2         CONV_FLASH_C20_ND+ CONV_N117524
+  CONV_FLASH_C20_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C20_M3         CONV_FLASH_C20_ND- CONV_FLASH_C20_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C62_M4         CONV_FLASH_C62_ND+ CONV_FLASH_C62_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C62_M5         CONV_FLASH_C62_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C62_M6         Q62 CONV_FLASH_C62_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C62_M7         Q62 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C62_M1         CONV_FLASH_C62_ND- N117007 CONV_FLASH_C62_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C62_M2         CONV_FLASH_C62_ND+ CONV_N119883
+  CONV_FLASH_C62_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C62_M3         CONV_FLASH_C62_ND- CONV_FLASH_C62_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C57_M4         CONV_FLASH_C57_ND+ CONV_FLASH_C57_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C57_M5         CONV_FLASH_C57_NDBIAS N117027 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
M_CONV_FLASH_C57_M6         Q57 CONV_FLASH_C57_ND+ N116990 N116990 CMOSP  
+ L=.2u  
+ W=.8u         
M_CONV_FLASH_C57_M7         Q57 N117027 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C57_M1         CONV_FLASH_C57_ND- N117007 CONV_FLASH_C57_NDBIAS 0
+  CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C57_M2         CONV_FLASH_C57_ND+ CONV_N119893
+  CONV_FLASH_C57_NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
M_CONV_FLASH_C57_M3         CONV_FLASH_C57_ND- CONV_FLASH_C57_ND- N116990
+  N116990 CMOSP  
+ L=.2u  
+ W=.6u         
R_CONV_1R-DIV_R42         CONV_N117534 CONV_N117532  10k  
R_CONV_1R-DIV_R15         CONV_N117490 CONV_N117488  10k  
R_CONV_1R-DIV_R55         CONV_N117558 CONV_N117556  10k  
R_CONV_1R-DIV_R63         CONV_1R-DIV_N02264 CONV_N117580  5k  
R_CONV_1R-DIV_R29         CONV_N117510 CONV_N117508  10k  
R_CONV_1R-DIV_R68         CONV_N117564 CONV_1R-DIV_N17274  5k  
R_CONV_1R-DIV_R43         CONV_N117536 CONV_N117534  10k  
R_CONV_1R-DIV_R56         CONV_N117560 CONV_N117558  10k  
R_CONV_1R-DIV_R30         CONV_N117512 CONV_N117510  10k  
R_CONV_1R-DIV_R16         CONV_N117492 CONV_N117490  10k  
R_CONV_1R-DIV_R70         CONV_1R-DIV_N169051 CONV_N117582  5k  
R_CONV_1R-DIV_R8         CONV_1R-DIV_R56 CONV_1R-DIV_R57  10k  
R_CONV_1R-DIV_R1         CONV_1R-DIV_R63 N117050  5k  
R_CONV_1R-DIV_R64         CONV_N117568 CONV_N117564  10k  
R_CONV_1R-DIV_R44         CONV_N117538 CONV_N117536  10k  
R_CONV_1R-DIV_R57         CONV_N117562 CONV_N117560  10k  
R_CONV_1R-DIV_R31         CONV_N117514 CONV_N117512  10k  
R_CONV_1R-DIV_R17         CONV_N117494 CONV_N117492  10k  
R_CONV_1R-DIV_R65         CONV_N117566 CONV_N117568  10k  
R_CONV_1R-DIV_R2         CONV_1R-DIV_R62 CONV_1R-DIV_R63  10k  
R_CONV_1R-DIV_R45         CONV_N117540 CONV_N117538  10k  
R_CONV_1R-DIV_R58         CONV_1R-DIV_N02264 CONV_N117562  5k  
R_CONV_1R-DIV_R18         CONV_N117496 CONV_N117494  10k  
R_CONV_1R-DIV_R32         CONV_N117516 CONV_N117514  10k  
R_CONV_1R-DIV_R66         CONV_N117574 CONV_N117566  10k  
R_CONV_1R-DIV_R9         CONV_1R-DIV_R55 CONV_1R-DIV_R56  10k  
R_CONV_1R-DIV_R46         CONV_N117542 CONV_N117540  10k  
R_CONV_1R-DIV_R3         CONV_1R-DIV_R61 CONV_1R-DIV_R62  10k  
R_CONV_1R-DIV_R19         CONV_N117498 CONV_N117496  10k  
R_CONV_1R-DIV_R33         CONV_N117518 CONV_N117516  10k  
R_CONV_1R-DIV_R67         CONV_N117572 CONV_N117574  10k  
R_CONV_1R-DIV_R47         CONV_N117544 CONV_N117542  10k  
R_CONV_1R-DIV_R20         CONV_N117500 CONV_N117498  10k  
R_CONV_1R-DIV_R34         CONV_N117520 CONV_N117518  10k  
R_CONV_1R-DIV_R69         CONV_N117582 CONV_1R-DIV_N17274  5k  
R_CONV_1R-DIV_R10         CONV_1R-DIV_R54 CONV_1R-DIV_R55  10k  
R_CONV_1R-DIV_R48         CONV_1R-DIV_N03146 CONV_N117544  5k  
R_CONV_1R-DIV_R21         CONV_1R-DIV_R50 CONV_N117500  10k  
R_CONV_1R-DIV_R4         CONV_1R-DIV_R60 CONV_1R-DIV_R61  10k  
R_CONV_1R-DIV_R35         CONV_N117522 CONV_N117520  10k  
R_CONV_1R-DIV_R49         CONV_N117546 CONV_1R-DIV_N03539  5k  
R_CONV_1R-DIV_R37         CONV_N117524 CONV_1R-DIV_N03539  5k  
R_CONV_1R-DIV_R22         CONV_1R-DIV_R51 CONV_1R-DIV_R50  10k  
R_CONV_1R-DIV_R50         CONV_N117548 CONV_N117546  10k  
R_CONV_1R-DIV_R36         CONV_1R-DIV_N03146 CONV_N117522  5k  
R_CONV_1R-DIV_R5         CONV_1R-DIV_R59 CONV_1R-DIV_R60  10k  
R_CONV_1R-DIV_R38         CONV_N117526 CONV_N117524  10k  
R_CONV_1R-DIV_R51         CONV_N117550 CONV_N117548  10k  
R_CONV_1R-DIV_R23         CONV_1R-DIV_R52 CONV_1R-DIV_R51  10k  
R_CONV_1R-DIV_R11         CONV_1R-DIV_R53 CONV_1R-DIV_R54  10k  
R_CONV_1R-DIV_R59         CONV_N117570 CONV_N117572  10k  
R_CONV_1R-DIV_R25         CONV_N117502 CONV_1R-DIV_N03082  5k  
R_CONV_1R-DIV_R39         CONV_N117528 CONV_N117526  10k  
R_CONV_1R-DIV_R24         CONV_1R-DIV_N03019 CONV_1R-DIV_R52  5k  
R_CONV_1R-DIV_R26         CONV_N117504 CONV_N117502  10k  
R_CONV_1R-DIV_R52         CONV_N117552 CONV_N117550  10k  
R_CONV_1R-DIV_R60         CONV_N117576 CONV_N117570  10k  
R_CONV_1R-DIV_R6         CONV_1R-DIV_R58 CONV_1R-DIV_R59  10k  
R_CONV_1R-DIV_R27         CONV_N117506 CONV_N117504  10k  
R_CONV_1R-DIV_R61         CONV_N117578 CONV_N117576  10k  
R_CONV_1R-DIV_R40         CONV_N117530 CONV_N117528  10k  
R_CONV_1R-DIV_R53         CONV_N117554 CONV_N117552  10k  
R_CONV_1R-DIV_R13         CONV_N117486 CONV_1R-DIV_N03082  5k  
V_CONV_1R-DIV_V1         CONV_1R-DIV_N169051 0 200mV
R_CONV_1R-DIV_R12         CONV_1R-DIV_N03019 CONV_1R-DIV_R53  5k  
R_CONV_1R-DIV_R41         CONV_N117532 CONV_N117530  10k  
R_CONV_1R-DIV_R54         CONV_N117556 CONV_N117554  10k  
R_CONV_1R-DIV_R14         CONV_N117488 CONV_N117486  10k  
R_CONV_1R-DIV_R62         CONV_N117580 CONV_N117578  10k  
R_CONV_1R-DIV_R28         CONV_N117508 CONV_N117506  10k  
R_CONV_1R-DIV_R7         CONV_1R-DIV_R57 CONV_1R-DIV_R58  10k  
R_CONV_2R-DIV_R42         CONV_2R-DIV_R25 CONV_2R-DIV_R24  10k  
R_CONV_2R-DIV_R15         CONV_2R-DIV_R44 CONV_2R-DIV_R43  10k  
R_CONV_2R-DIV_R55         CONV_2R-DIV_R13 CONV_2R-DIV_R14  10k  
R_CONV_2R-DIV_R63         CONV_2R-DIV_N02264 CONV_2R-DIV_R10  5k  
R_CONV_2R-DIV_R29         CONV_2R-DIV_R37 CONV_2R-DIV_R38  10k  
R_CONV_2R-DIV_R68         CONV_2R-DIV_R2 CONV_2R-DIV_N17274  5k  
R_CONV_2R-DIV_R43         CONV_2R-DIV_R26 CONV_2R-DIV_R25  10k  
R_CONV_2R-DIV_R56         CONV_2R-DIV_R12 CONV_2R-DIV_R13  10k  
R_CONV_2R-DIV_R30         CONV_2R-DIV_R36 CONV_2R-DIV_R37  10k  
R_CONV_2R-DIV_R16         CONV_2R-DIV_R45 CONV_2R-DIV_R44  10k  
R_CONV_2R-DIV_R70         CONV_2R-DIV_N169051 CONV_2R-DIV_R1  5k  
R_CONV_2R-DIV_R8         CONV_N119895 CONV_N119893  10k  
R_CONV_2R-DIV_R1         CONV_N119881 N117050  5k  
R_CONV_2R-DIV_R64         CONV_2R-DIV_R3 CONV_2R-DIV_R2  10k  
R_CONV_2R-DIV_R44         CONV_2R-DIV_R27 CONV_2R-DIV_R26  10k  
R_CONV_2R-DIV_R57         CONV_2R-DIV_R11 CONV_2R-DIV_R12  10k  
R_CONV_2R-DIV_R31         CONV_2R-DIV_R35 CONV_2R-DIV_R36  10k  
R_CONV_2R-DIV_R17         CONV_2R-DIV_R46 CONV_2R-DIV_R45  10k  
R_CONV_2R-DIV_R65         CONV_2R-DIV_R4 CONV_2R-DIV_R3  10k  
R_CONV_2R-DIV_R2         CONV_N119883 CONV_N119881  10k  
R_CONV_2R-DIV_R45         CONV_2R-DIV_R28 CONV_2R-DIV_R27  10k  
R_CONV_2R-DIV_R58         CONV_2R-DIV_N02264 CONV_2R-DIV_R11  5k  
R_CONV_2R-DIV_R18         CONV_2R-DIV_R47 CONV_2R-DIV_R46  10k  
R_CONV_2R-DIV_R32         CONV_2R-DIV_R34 CONV_2R-DIV_R35  10k  
R_CONV_2R-DIV_R66         CONV_2R-DIV_R5 CONV_2R-DIV_R4  10k  
R_CONV_2R-DIV_R9         CONV_N119897 CONV_N119895  10k  
R_CONV_2R-DIV_R46         CONV_2R-DIV_R29 CONV_2R-DIV_R28  10k  
R_CONV_2R-DIV_R3         CONV_N119885 CONV_N119883  10k  
R_CONV_2R-DIV_R19         CONV_2R-DIV_R48 CONV_2R-DIV_R47  10k  
R_CONV_2R-DIV_R33         CONV_2R-DIV_R33 CONV_2R-DIV_R34  10k  
R_CONV_2R-DIV_R67         CONV_2R-DIV_R6 CONV_2R-DIV_R5  10k  
R_CONV_2R-DIV_R47         CONV_2R-DIV_R30 CONV_2R-DIV_R29  10k  
R_CONV_2R-DIV_R20         CONV_2R-DIV_R49 CONV_2R-DIV_R48  10k  
R_CONV_2R-DIV_R34         CONV_2R-DIV_R32 CONV_2R-DIV_R33  10k  
R_CONV_2R-DIV_R69         CONV_2R-DIV_R1 CONV_2R-DIV_N17274  5k  
R_CONV_2R-DIV_R10         CONV_N119899 CONV_N119897  10k  
R_CONV_2R-DIV_R48         CONV_2R-DIV_N03146 CONV_2R-DIV_R30  5k  
R_CONV_2R-DIV_R21         CONV_N119903 CONV_2R-DIV_R49  10k  
R_CONV_2R-DIV_R4         CONV_N119887 CONV_N119885  10k  
R_CONV_2R-DIV_R35         CONV_2R-DIV_R31 CONV_2R-DIV_R32  10k  
R_CONV_2R-DIV_R49         CONV_2R-DIV_R19 CONV_2R-DIV_N03539  5k  
R_CONV_2R-DIV_R37         CONV_2R-DIV_R20 CONV_2R-DIV_N03539  5k  
R_CONV_2R-DIV_R22         CONV_N119905 CONV_N119903  10k  
R_CONV_2R-DIV_R50         CONV_2R-DIV_R18 CONV_2R-DIV_R19  10k  
R_CONV_2R-DIV_R36         CONV_2R-DIV_N03146 CONV_2R-DIV_R31  5k  
R_CONV_2R-DIV_R5         CONV_N119889 CONV_N119887  10k  
R_CONV_2R-DIV_R38         CONV_2R-DIV_R21 CONV_2R-DIV_R20  10k  
R_CONV_2R-DIV_R51         CONV_2R-DIV_R17 CONV_2R-DIV_R18  10k  
R_CONV_2R-DIV_R23         CONV_N119907 CONV_N119905  10k  
R_CONV_2R-DIV_R11         CONV_N119901 CONV_N119899  10k  
R_CONV_2R-DIV_R59         CONV_2R-DIV_R7 CONV_2R-DIV_R6  10k  
R_CONV_2R-DIV_R25         CONV_2R-DIV_R41 CONV_2R-DIV_N03082  5k  
R_CONV_2R-DIV_R39         CONV_2R-DIV_R22 CONV_2R-DIV_R21  10k  
R_CONV_2R-DIV_R24         CONV_2R-DIV_N03019 CONV_N119907  5k  
R_CONV_2R-DIV_R26         CONV_2R-DIV_R40 CONV_2R-DIV_R41  10k  
R_CONV_2R-DIV_R52         CONV_2R-DIV_R16 CONV_2R-DIV_R17  10k  
R_CONV_2R-DIV_R60         CONV_2R-DIV_R8 CONV_2R-DIV_R7  10k  
R_CONV_2R-DIV_R6         CONV_N119891 CONV_N119889  10k  
R_CONV_2R-DIV_R27         CONV_2R-DIV_R39 CONV_2R-DIV_R40  10k  
R_CONV_2R-DIV_R61         CONV_2R-DIV_R9 CONV_2R-DIV_R8  10k  
R_CONV_2R-DIV_R40         CONV_2R-DIV_R23 CONV_2R-DIV_R22  10k  
R_CONV_2R-DIV_R53         CONV_2R-DIV_R15 CONV_2R-DIV_R16  10k  
R_CONV_2R-DIV_R13         CONV_2R-DIV_R42 CONV_2R-DIV_N03082  5k  
V_CONV_2R-DIV_V1         CONV_2R-DIV_N169051 0 200mV
R_CONV_2R-DIV_R12         CONV_2R-DIV_N03019 CONV_N119901  5k  
R_CONV_2R-DIV_R41         CONV_2R-DIV_R24 CONV_2R-DIV_R23  10k  
R_CONV_2R-DIV_R54         CONV_2R-DIV_R14 CONV_2R-DIV_R15  10k  
R_CONV_2R-DIV_R14         CONV_2R-DIV_R43 CONV_2R-DIV_R42  10k  
R_CONV_2R-DIV_R62         CONV_2R-DIV_R10 CONV_2R-DIV_R9  10k  
R_CONV_2R-DIV_R28         CONV_2R-DIV_R38 CONV_2R-DIV_R39  10k  
R_CONV_2R-DIV_R7         CONV_N119893 CONV_N119891  10k  
R_R9         N-4SB N116990  100k  
V_VBIAS         N117027 0 .33
R_R10         N-3SB N116990  100k  
R_R11         N-2SB N116990  100k  
V_VDD         N116990 0 3.3
V_VREF         N117050 0 3.035
R_R12         N-LSB N116990  100k  
V_VA         N117007 0 3
R_R1         MSB N116990  100k  
R_R2         5SB N116990  100k  
R_R3         4SB N116990  100k  
R_R4         3SB N116990  100k  
R_R5         2SB N116990  100k  