LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY SCHEMATIC1 IS 

END SCHEMATIC1;



ARCHITECTURE STRUCTURE OF SCHEMATIC1 IS

-- COMPONENTS

-- SIGNALS

SIGNAL \0\ : std_logic;
SIGNAL GND_0 : std_logic;

-- INSTANCE ATTRIBUTES



-- GATE INSTANCES

BEGIN
GND_0<=\0\;
GND_0<=\0\;
END STRUCTURE;

