
**** 04/17/10 16:10:21 ******* PSpice 16.0.0 (July 2006) ****** ID# 0 ********

 ** Profile: "TEST-transient"  [ D:\Documents\TESIS\fiocs\Design\I-COMPARADOR-02\OrCAD\i-comparador-01-pspicefiles\test\transient.sim


 ****     CIRCUIT DESCRIPTION


******************************************************************************




** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:\Documents\TESIS\fiocs\Design\I-COMPARADOR-02\OrCAD\I-COMPARADOR-01-PSpiceFiles/i-comparador-01.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.0\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 

.STEP V_VIN LIST 0.5 0.99 1 1.01 1.5
.TRAN  0 150n 0 10p 
.PROBE V(*) I(*) 

*.INC "..\TEST.net" 



**** INCLUDING TEST.net ****
* source I-COMPARADOR-01

M_M2         ND+ IN+ NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
V_VREF         IN+ N398131 1
M_M3         ND- ND- N39211 N39211 CMOSP  
+ L=.2u  
+ W=.6u         
M_M4         ND+ ND- N39211 N39211 CMOSP  
+ L=.2u  
+ W=.6u         
M_M5         NDBIAS VBIAS 0 0 CMOSN  
+ L=.2u  
+ W=.6u         
C_C1         0 N749310  1n  
V_VQ+         N398131 0 .2
M_U2_M5         N75001 NOUT N39211 N39211 CMOSP  
+ L=.18u  
+ W=.2u         
M_U2_M6         N75001 NOUT 0 0 CMOSN  
+ L=.18u  
+ W=.18u         
M_M6         NOUT ND+ N39211 N39211 CMOSP  
+ L=.2u  
+ W=.8u         
V_VBIAS         VBIAS 0 .33
M_M7         NOUT VBIAS 0 0 CMOSN  
+ L=.2u  
+ W=.4u         
V_VQ-         N43113 0 .2
V_VIN         IN- N43113 1.5
R_R1         N75001 N749310  500k  
M_M1         ND- IN- NDBIAS 0 CMOSN  
+ L=.2u  
+ W=.4u         
V_VDD         N39211 0 3.3

I_I1         ND+ 0 DC 0Adc AC 0Aac
+PULSE 0 4m 2n 50p 1.55n 100p 0


.END