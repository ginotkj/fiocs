** Profile: "PRUEBA-transient"  [ D:\Documents\TESIS\fiocs\Design\I-FLASH-01\OrCAD\I-FLASH-6BITS\i-flash-6bits-PSpiceFiles\PRUEBA\transient.sim ] 

** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../i-flash-6bits-pspicefiles/i-flash-6bits.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.0\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 15n 0 1p 
.OPTIONS NODE
.OPTIONS ITL1= 300
.OPTIONS ITL2= 100
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\PRUEBA.net" 


.END
