I_I1         N44303 0 DC 0Adc AC 0Aac 
 +EXP 0 4m 2n 30p 2.2n 500p
.PROBE/CSDF I(+EXP 0 4m 2n 30p 2.2n 500p)
.PROBE/CSDF ID(M_M2) IB(M_M2) IS(M_M2) IG(M_M2)
.PROBE/CSDF ID(M_M1) IB(M_M1) IS(M_M1) IG(M_M1)
.PROBE/CSDF ID(M_M5) IB(M_M5) IS(M_M5) IG(M_M5)
.END