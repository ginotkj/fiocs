-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Sunday, April 12, 2009 20:05:17 Argentina Standard Time

