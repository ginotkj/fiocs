****************************
*MODEL OF TANSISTORS    *
****************************
.MODEL NMOS NMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 3.12E-8
+XJ      = 3E-7           NCH     = 7.5E16         VTH0    = 0.5525942
+K1      = 0.9684018      K2      = -0.087558      K3      = 4.6086605
+K3B     = -2.0128057     W0      = 6.714563E-7    NLX     = 1.217197E-8
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.5293567      DVT1    = 0.4432139      DVT2    = -0.5
+U0      = 649.4788739    UA      = 1.313648E-9    UB      = 2.836687E-18
+UC      = 2.458363E-11   VSAT    = 1.170587E5     A0      = 0.6528338
+AGS     = 0.1136675      B0      = 1.489912E-6    B1      = 5E-6
+KETA    = -8.095926E-3   A1      = 0              A2      = 1
+RDSW    = 3E3            PRWG    = -5.073199E-4   PRWB    = -0.0618845
+WR      = 1              WINT    = 7.755726E-7    LINT    = 1.819685E-7
+XL      = 0              XW      = 0              DWG     = -2.496315E-8
+DWB     = 1.669565E-8    VOFF    = -0.0731456     NFACTOR = 0.567383
+CIT     = 0              CDSC    = 7.627884E-6    CDSCD   = 8.475154E-6
+CDSCB   = 4.691294E-5    ETA0    = -0.6101195     ETAB    = -0.300202
+DSUB    = 0.8799726      PCLM    = 1.8481182      PDIBLC1 = 8.801319E-3
+PDIBLC2 = 1.58414E-3     PDIBLCB = -0.1           DROUT   = 0.0681381
+PSCBE1  = 6.290635E9     PSCBE2  = 1.441641E-9    PVAG    = 0.91451
+DELTA   = 0.01           RSH     = 52.7           MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 1.75E-10       CGSO    = 1.75E-10       CGBO    = 1E-9
+CJ      = 2.737552E-4    PB      = 0.99           MJ      = 0.5481931
+CJSW    = 1.359277E-10   PBSW    = 0.99           MJSW    = 0.1
+CJSWG   = 6.4E-11        PBSWG   = 0.99           MJSWG   = 0.1
+CF      = 0               )
*
*.MODEL Dpdiff D RS=1
.MODEL PMOS PMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 3.12E-8
+XJ      = 3E-7           NCH     = 2.4E16         VTH0    = -0.8476404
+K1      = 0.4513608      K2      = 2.379699E-5    K3      = 13.3278347
+K3B     = -2.2238332     W0      = 9.577236E-7    NLX     = 1E-6
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.4907854      DVT1    = 0.665622       DVT2    = -0.0372218
+U0      = 236.8923827    UA      = 3.833306E-9    UB      = 1.487688E-21
+UC      = -1.08562E-10   VSAT    = 2E5            A0      = 0.4205945
+AGS     = 0.2140979      B0      = 6.620808E-6    B1      = 5E-6
+KETA    = 5.754484E-3    A1      = 0              A2      = 0.364
+RDSW    = 3E3            PRWG    = 0.2425124      PRWB    = -0.2108462
+WR      = 1              WINT    = 7.565065E-7    LINT    = 3.218813E-8
+XL      = 0              XW      = 0              DWG     = -2.13917E-8
+DWB     = 3.857544E-8    VOFF    = -0.0877184     NFACTOR = 0.2508342
+CIT     = 0              CDSC    = 2.924806E-5    CDSCD   = 1.497572E-4
+CDSCB   = 1.091488E-4    ETA0    = 0.26103        ETAB    = -8.148244E-4
+DSUB    = 0.2873         PCLM    = 1.120595E-10   PDIBLC1 = 4.502478E-4
+PDIBLC2 = 1.090076E-3    PDIBLCB = -1E-3          DROUT   = 9.243538E-4
+PSCBE1  = 3.500883E9     PSCBE2  = 5.252383E-10   PVAG    = 15
+DELTA   = 0.01           RSH     = 76             MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.1E-10        CGSO    = 2.1E-10        CGBO    = 1E-9
+CJ      = 3.085988E-4    PB      = 0.8            MJ      = 0.4394529
+CJSW    = 1.58319E-10    PBSW    = 0.9882954      MJSW    = 0.1003165
+CJSWG   = 3.9E-11        PBSWG   = 0.9882954      MJSWG   = 0.1003165
+CF      = 0               )
**
