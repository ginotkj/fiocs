** Profile: "S-NAND-3-bias1"  [ D:\Documents\TESIS\TRUNK\Design\I-FFD-01\i-ffd-01-pspicefiles\s-nand-3\bias1.sim ] 

** Creating circuit file "bias1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_10.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\S-NAND-3.net" 


.END
