I_I1         N48205 0 DC 0Adc AC 0Aac 
 +EXP 0 4m 2n 30p 2.2n 500p
.PROBE/CSDF I(+EXP 0 4m 2n 30p 2.2n 500p)
.PROBE/CSDF ID(M_M9) IB(M_M9) IS(M_M9) IG(M_M9)
.PROBE/CSDF ID(M_M2) IB(M_M2) IS(M_M2) IG(M_M2)
.PROBE/CSDF ID(M_M4) IB(M_M4) IS(M_M4) IG(M_M4)
.END