** Profile: "Tech-1.6um-Tech-1.6um"  [ C:\Documents and Settings\fjferre1\My Documents\NOBACKUP\Tesis\Repo\Design\E-OPAMP-001\E-OPAMP-001-PSpiceFiles\Tech-1.6um\Tech-1.6um.sim ] 

** Creating circuit file "Tech-1.6um.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../e-opamp-001-pspicefiles/e-opamp-001.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.2\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OP
.SAVEBIAS "./bias_tech-1_6.txt" OP 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Tech-1.6um.net" 


.END
