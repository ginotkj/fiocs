**** 05/12/10 18:10:37 ******* PSpice 16.0.0 (July 2006) ****** ID# 0 ********

 ** Profile: "DOBLE-NEG-PRUEBA"  [ D:\Documents\TESIS\fiocs\Design\I-COMPARADOR-01\OrCAD\i-comparador-01-pspicefiles\doble-neg\prueba

 ****     CIRCUIT DESCRIPTION
******************************************************************************

* Local Libraries :
.LIB "D:\Documents\TESIS\fiocs\Design\I-COMPARADOR-01\OrCAD\i-comparador-01-pspicefiles\i-comparador-01.lib" 
.lib "nom.lib" 

*Analysis directives: 
.STEP V_VIN LIST -10m -5m 5m 10m
.TRAN  0 100n 0 0 
.PROBE V(*) I(*) 

**** INCLUDING DOBLE-NEG.net ****
* source I-COMPARADOR-01

V_VIN         VINNEG N652820 0
M_M1         NDNEG VINNEG NDBIAS 0 CMOSN  
+ L=10u  
+ W=265u         
M_M2         NDPOS VINPOS NDBIAS 0 CMOSN  
+ L=10u  
+ W=265u         
V_VDD         N64870 0 3.3
M_M3         NDNEG NDNEG N64870 N64870 CMOSP  
+ L=10u  
+ W=200u         
V_VBIAS         VBIAS 0 1
M_M12         NDOUT NDPOS N64870 N64870 CMOSP  
+ L=10u  
+ W=1120u         
V_VQ2         N1312720 0 1.320
M_M4         NDPOS NDNEG N64870 N64870 CMOSP  
+ L=10u  
+ W=200u         
M_M13         NDOUT VBIAS 0 0 CMOSN  
+ L=15u  
+ W=220u         
M_M5         NDBIAS VBIAS 0 0 CMOSN  
+ L=12.5u  
+ W=65u         
V_VQ1         N652820 0 1.320
V_VREF         VINPOS N1312720 0

I_INYECCION	0 NDOUT DC 0Adc AC 0Aac
+EXP 0 2m 2n 80p 5.5n 1n

.END