** Profile: "SCHEMATIC1-bias"  [ D:\DOCUMENTS\TESIS\TRUNK\DESIGN\I-COMPARADOR-01\i-comparador-01-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../i-comparador-01-pspicefiles/i-comparador-01.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\OrCAD 16\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
