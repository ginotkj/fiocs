**** 05/12/10 18:10:37 ******* PSpice 16.0.0 (July 2006) ****** ID# 0 ********

 ** Profile: "DOBLE-NEG-PRUEBA"  [ D:\Documents\TESIS\fiocs\Design\I-COMPARADOR-01\OrCAD\i-comparador-01-pspicefiles\doble-neg\prueba

 ****     CIRCUIT DESCRIPTION
******************************************************************************

* Local Libraries :
.LIB "D:\Documents\TESIS\fiocs\Design\I-COMPARADOR-01\OrCAD\i-comparador-01-pspicefiles\i-comparador-01.lib" 
.lib "nom.lib" 

*Analysis directives: 
.STEP V_VIN LIST 1.05 1.055 1.065 1.07
.TRAN  0 100n 0 0 
.PROBE V(*) I(*) 

**** INCLUDING DOBLE-NEG.net ****
* source I-COMPARADOR-01

M_M1         NDNEG VINNEG NDBIAS 0 CMOSN  
+ L=20u  
+ W=89u         
M_M2         NDPOS VINPOS NDBIAS 0 CMOSN  
+ L=20u  
+ W=89u         
V_VDD         N64870 0 3.3
M_M3         NDNEG NDNEG N64870 N64870 CMOSP  
+ L=25u  
+ W=37u         
V_VBIAS         VBIAS 0 .52
M_M12         NDOUT NDPOS N64870 N64870 CMOSP  
+ L=15u  
+ W=1097u         
M_M4         NDPOS NDNEG N64870 N64870 CMOSP  
+ L=25u  
+ W=37u         
M_M13         NDOUT VBIAS 0 0 CMOSN  
+ L=15u  
+ W=375u         
M_M5         NDBIAS VBIAS 0 0 CMOSN  
+ L=20u  
+ W=20u         
V_VIN         VINNEG 0 1.063    
V_VREF         VINPOS 0 1.063              


I_INYECCION	0 NDNEG DC 0Adc AC 0Aac
+EXP 0 2m 2n 80p 5.5n 1n

.END