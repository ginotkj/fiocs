I_I1         N73485 0 DC 0Adc AC 0Aac 
 +EXP 0 4m 2n 30p 2.2n 500p
.PROBE/CSDF I(+EXP 0 4m 2n 30p 2.2n 500p)
.PROBE/CSDF ID(M_M12) IB(M_M12) IS(M_M12) IG(M_M12)
.PROBE/CSDF ID(M_M11) IB(M_M11) IS(M_M11) IG(M_M11)
.END