** Profile: "SCHEMATIC1-bode"  [ D:\DOCUMENTS\TESIS\TRUNK\DESIGN\I-PBFILTER-01\I-PBFILTER-01-PSpiceFiles\SCHEMATIC1\bode.sim ] 

** Creating circuit file "bode.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../i-pbfilter-01-pspicefiles/i-pbfilter-01.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.2\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 1 100G
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
