** Profile: "SCHEMATIC1-ac"  [ D:\DOCUMENTS\TESIS\TRUNK\DESIGN\I-OPAMPB-01\I-OPAMPB-01-PSpiceFiles\SCHEMATIC1\ac.sim ] 

** Creating circuit file "ac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../i-opampb-01-pspicefiles/i-opampb-01.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.2\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 10 10 1M
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
