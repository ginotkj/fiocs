*******************************
* Begin .SUBCKT model         *
* spice-sdb ver 4.28.2007     *
*******************************
.SUBCKT 2nand1 1 6 2 4 5 
*vvvvvvvv  Included SPICE model from ../model/pmos.model vvvvvvvv
.model mos_p PMOS(LEVEL=3 PHI=0.600000 TOX=2.1200E-08 XJ=0.200000U 
+  TPG=-1 VTO=-0.9056 DELTA=1.5200E+00 LD=2.2000E-08 KP=2.9352E-05
+  UO=180.2 THETA=1.2480E-01 RSH=1.0470E+02 GAMMA=0.4863
+  NSUB=1.8900E+16 NFS=3.46E+12 VMAX=3.7320E+05 ETA=1.6410E-01
+  KAPPA=9.6940E+00 CGDO=5.3752E-11 CGSO=5.3752E-11
+  CGBO=3.3650E-10 CJ=4.8447E-04 MJ=0.5027 CJSW=1.6457E-10
+  MJSW=0.217168 PB=0.850000)
*^^^^^^^^  End of included SPICE model from ../model/pmos.model ^^^^^^^^
*
*==============  Begin SPICE netlist of main design ============
M4 1 5 6 6 pmos4  l=1u w=10u
M3 1 4 6 6 pmos4  l=1u w=10u
M2 3 5 2 2 nmos4  l=3u w=1u
M1 1 4 3 2 nmos4  l=3u w=1u
.ends 2nand1
*******************************
