I_I1         N55353 0 DC 0Adc AC 0Aac 
 +EXP 0 4m 2n 30p 2.2n 500p
.PROBE/CSDF I(+EXP 0 4m 2n 30p 2.2n 500p)
.PROBE/CSDF ID(M_M10) IB(M_M10) IS(M_M10) IG(M_M10)
.PROBE/CSDF ID(M_M9) IB(M_M9) IS(M_M9) IG(M_M9)
.PROBE/CSDF ID(M_M8) IB(M_M8) IS(M_M8) IG(M_M8)
.PROBE/CSDF ID(M_M7) IB(M_M7) IS(M_M7) IG(M_M7)
.END